// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 24 2015 00:15:54

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSync,
    SDATA,
    SCLK1,
    Pixel,
    HSync,
    nCS2,
    SCLK2,
    Clock12MHz,
    nCS1);

    output VSync;
    input SDATA;
    output SCLK1;
    output Pixel;
    output HSync;
    output nCS2;
    output SCLK2;
    input Clock12MHz;
    output nCS1;

    wire N__16513;
    wire N__16512;
    wire N__16511;
    wire N__16502;
    wire N__16501;
    wire N__16500;
    wire N__16493;
    wire N__16492;
    wire N__16491;
    wire N__16484;
    wire N__16483;
    wire N__16482;
    wire N__16475;
    wire N__16474;
    wire N__16473;
    wire N__16466;
    wire N__16465;
    wire N__16464;
    wire N__16457;
    wire N__16456;
    wire N__16455;
    wire N__16448;
    wire N__16447;
    wire N__16446;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16403;
    wire N__16402;
    wire N__16401;
    wire N__16398;
    wire N__16397;
    wire N__16396;
    wire N__16395;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16384;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16364;
    wire N__16361;
    wire N__16356;
    wire N__16355;
    wire N__16352;
    wire N__16349;
    wire N__16348;
    wire N__16343;
    wire N__16340;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16319;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16303;
    wire N__16294;
    wire N__16291;
    wire N__16286;
    wire N__16281;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16236;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16221;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16209;
    wire N__16208;
    wire N__16207;
    wire N__16204;
    wire N__16203;
    wire N__16202;
    wire N__16201;
    wire N__16200;
    wire N__16199;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16191;
    wire N__16190;
    wire N__16187;
    wire N__16186;
    wire N__16185;
    wire N__16184;
    wire N__16183;
    wire N__16180;
    wire N__16173;
    wire N__16166;
    wire N__16157;
    wire N__16156;
    wire N__16155;
    wire N__16154;
    wire N__16153;
    wire N__16152;
    wire N__16151;
    wire N__16148;
    wire N__16139;
    wire N__16138;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16112;
    wire N__16107;
    wire N__16104;
    wire N__16099;
    wire N__16096;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16074;
    wire N__16073;
    wire N__16072;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16029;
    wire N__16028;
    wire N__16025;
    wire N__16024;
    wire N__16023;
    wire N__16022;
    wire N__16021;
    wire N__16020;
    wire N__16019;
    wire N__16018;
    wire N__16017;
    wire N__16016;
    wire N__16015;
    wire N__16014;
    wire N__16013;
    wire N__16012;
    wire N__16011;
    wire N__16010;
    wire N__16009;
    wire N__16008;
    wire N__16007;
    wire N__16006;
    wire N__16005;
    wire N__16004;
    wire N__16003;
    wire N__16002;
    wire N__16001;
    wire N__16000;
    wire N__15999;
    wire N__15998;
    wire N__15997;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15985;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15975;
    wire N__15972;
    wire N__15965;
    wire N__15962;
    wire N__15955;
    wire N__15950;
    wire N__15945;
    wire N__15936;
    wire N__15927;
    wire N__15920;
    wire N__15919;
    wire N__15918;
    wire N__15917;
    wire N__15912;
    wire N__15905;
    wire N__15898;
    wire N__15891;
    wire N__15888;
    wire N__15875;
    wire N__15870;
    wire N__15869;
    wire N__15868;
    wire N__15867;
    wire N__15866;
    wire N__15863;
    wire N__15862;
    wire N__15861;
    wire N__15854;
    wire N__15851;
    wire N__15844;
    wire N__15841;
    wire N__15828;
    wire N__15817;
    wire N__15816;
    wire N__15815;
    wire N__15814;
    wire N__15813;
    wire N__15812;
    wire N__15809;
    wire N__15808;
    wire N__15807;
    wire N__15806;
    wire N__15805;
    wire N__15804;
    wire N__15803;
    wire N__15800;
    wire N__15797;
    wire N__15796;
    wire N__15795;
    wire N__15794;
    wire N__15793;
    wire N__15792;
    wire N__15791;
    wire N__15790;
    wire N__15789;
    wire N__15784;
    wire N__15779;
    wire N__15776;
    wire N__15771;
    wire N__15770;
    wire N__15769;
    wire N__15762;
    wire N__15761;
    wire N__15760;
    wire N__15759;
    wire N__15758;
    wire N__15757;
    wire N__15756;
    wire N__15755;
    wire N__15754;
    wire N__15753;
    wire N__15748;
    wire N__15737;
    wire N__15734;
    wire N__15729;
    wire N__15728;
    wire N__15723;
    wire N__15718;
    wire N__15713;
    wire N__15710;
    wire N__15697;
    wire N__15696;
    wire N__15695;
    wire N__15694;
    wire N__15693;
    wire N__15692;
    wire N__15685;
    wire N__15684;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15664;
    wire N__15659;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15622;
    wire N__15619;
    wire N__15618;
    wire N__15617;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15609;
    wire N__15608;
    wire N__15605;
    wire N__15602;
    wire N__15595;
    wire N__15594;
    wire N__15593;
    wire N__15592;
    wire N__15591;
    wire N__15590;
    wire N__15589;
    wire N__15588;
    wire N__15587;
    wire N__15586;
    wire N__15585;
    wire N__15584;
    wire N__15581;
    wire N__15580;
    wire N__15579;
    wire N__15578;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15563;
    wire N__15560;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15545;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15521;
    wire N__15512;
    wire N__15505;
    wire N__15500;
    wire N__15499;
    wire N__15496;
    wire N__15493;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15475;
    wire N__15472;
    wire N__15467;
    wire N__15464;
    wire N__15457;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15429;
    wire N__15426;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15405;
    wire N__15404;
    wire N__15403;
    wire N__15402;
    wire N__15401;
    wire N__15400;
    wire N__15399;
    wire N__15398;
    wire N__15397;
    wire N__15396;
    wire N__15395;
    wire N__15394;
    wire N__15393;
    wire N__15390;
    wire N__15389;
    wire N__15386;
    wire N__15385;
    wire N__15384;
    wire N__15383;
    wire N__15382;
    wire N__15381;
    wire N__15380;
    wire N__15377;
    wire N__15376;
    wire N__15375;
    wire N__15368;
    wire N__15357;
    wire N__15356;
    wire N__15355;
    wire N__15354;
    wire N__15349;
    wire N__15338;
    wire N__15337;
    wire N__15336;
    wire N__15335;
    wire N__15334;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15326;
    wire N__15323;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15302;
    wire N__15301;
    wire N__15300;
    wire N__15299;
    wire N__15298;
    wire N__15297;
    wire N__15296;
    wire N__15295;
    wire N__15294;
    wire N__15289;
    wire N__15288;
    wire N__15287;
    wire N__15282;
    wire N__15277;
    wire N__15272;
    wire N__15269;
    wire N__15262;
    wire N__15259;
    wire N__15250;
    wire N__15249;
    wire N__15244;
    wire N__15241;
    wire N__15234;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15217;
    wire N__15214;
    wire N__15205;
    wire N__15200;
    wire N__15197;
    wire N__15190;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15148;
    wire N__15145;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15126;
    wire N__15121;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15102;
    wire N__15099;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15093;
    wire N__15090;
    wire N__15085;
    wire N__15082;
    wire N__15081;
    wire N__15078;
    wire N__15077;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15034;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15015;
    wire N__15014;
    wire N__15013;
    wire N__15012;
    wire N__15011;
    wire N__15010;
    wire N__15009;
    wire N__15008;
    wire N__15007;
    wire N__15004;
    wire N__15003;
    wire N__15000;
    wire N__14999;
    wire N__14996;
    wire N__14995;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14987;
    wire N__14986;
    wire N__14985;
    wire N__14984;
    wire N__14977;
    wire N__14976;
    wire N__14975;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14960;
    wire N__14955;
    wire N__14954;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14946;
    wire N__14943;
    wire N__14940;
    wire N__14935;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14920;
    wire N__14917;
    wire N__14914;
    wire N__14909;
    wire N__14904;
    wire N__14903;
    wire N__14902;
    wire N__14901;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14843;
    wire N__14836;
    wire N__14829;
    wire N__14822;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14778;
    wire N__14777;
    wire N__14776;
    wire N__14775;
    wire N__14774;
    wire N__14773;
    wire N__14770;
    wire N__14769;
    wire N__14768;
    wire N__14767;
    wire N__14766;
    wire N__14765;
    wire N__14762;
    wire N__14761;
    wire N__14760;
    wire N__14759;
    wire N__14758;
    wire N__14757;
    wire N__14754;
    wire N__14753;
    wire N__14752;
    wire N__14751;
    wire N__14750;
    wire N__14747;
    wire N__14746;
    wire N__14745;
    wire N__14744;
    wire N__14743;
    wire N__14742;
    wire N__14741;
    wire N__14738;
    wire N__14737;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14714;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14702;
    wire N__14695;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14676;
    wire N__14673;
    wire N__14666;
    wire N__14657;
    wire N__14652;
    wire N__14645;
    wire N__14642;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14634;
    wire N__14631;
    wire N__14630;
    wire N__14627;
    wire N__14622;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14599;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14582;
    wire N__14577;
    wire N__14574;
    wire N__14569;
    wire N__14564;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14458;
    wire N__14455;
    wire N__14452;
    wire N__14451;
    wire N__14450;
    wire N__14447;
    wire N__14446;
    wire N__14445;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14430;
    wire N__14427;
    wire N__14426;
    wire N__14425;
    wire N__14420;
    wire N__14415;
    wire N__14412;
    wire N__14407;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14388;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14361;
    wire N__14360;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14328;
    wire N__14327;
    wire N__14326;
    wire N__14325;
    wire N__14314;
    wire N__14311;
    wire N__14308;
    wire N__14307;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14278;
    wire N__14275;
    wire N__14272;
    wire N__14269;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14256;
    wire N__14255;
    wire N__14254;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14246;
    wire N__14245;
    wire N__14244;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14221;
    wire N__14218;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14206;
    wire N__14203;
    wire N__14196;
    wire N__14191;
    wire N__14184;
    wire N__14179;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14097;
    wire N__14094;
    wire N__14093;
    wire N__14090;
    wire N__14089;
    wire N__14086;
    wire N__14079;
    wire N__14074;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14062;
    wire N__14059;
    wire N__14058;
    wire N__14057;
    wire N__14054;
    wire N__14049;
    wire N__14048;
    wire N__14043;
    wire N__14040;
    wire N__14039;
    wire N__14038;
    wire N__14033;
    wire N__14032;
    wire N__14031;
    wire N__14030;
    wire N__14025;
    wire N__14022;
    wire N__14017;
    wire N__14014;
    wire N__14005;
    wire N__14004;
    wire N__14003;
    wire N__14000;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13911;
    wire N__13910;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13887;
    wire N__13886;
    wire N__13885;
    wire N__13882;
    wire N__13877;
    wire N__13876;
    wire N__13873;
    wire N__13872;
    wire N__13869;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13842;
    wire N__13839;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13749;
    wire N__13748;
    wire N__13741;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13719;
    wire N__13716;
    wire N__13715;
    wire N__13714;
    wire N__13713;
    wire N__13710;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13690;
    wire N__13689;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13663;
    wire N__13660;
    wire N__13659;
    wire N__13658;
    wire N__13657;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13645;
    wire N__13642;
    wire N__13633;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13618;
    wire N__13615;
    wire N__13612;
    wire N__13611;
    wire N__13608;
    wire N__13607;
    wire N__13604;
    wire N__13603;
    wire N__13600;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13564;
    wire N__13561;
    wire N__13552;
    wire N__13549;
    wire N__13546;
    wire N__13543;
    wire N__13542;
    wire N__13541;
    wire N__13540;
    wire N__13537;
    wire N__13536;
    wire N__13533;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13513;
    wire N__13510;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13495;
    wire N__13492;
    wire N__13489;
    wire N__13486;
    wire N__13483;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13471;
    wire N__13468;
    wire N__13465;
    wire N__13464;
    wire N__13461;
    wire N__13460;
    wire N__13459;
    wire N__13458;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13444;
    wire N__13441;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13423;
    wire N__13422;
    wire N__13419;
    wire N__13418;
    wire N__13417;
    wire N__13414;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13381;
    wire N__13378;
    wire N__13375;
    wire N__13372;
    wire N__13369;
    wire N__13366;
    wire N__13363;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13335;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13318;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13306;
    wire N__13305;
    wire N__13304;
    wire N__13303;
    wire N__13302;
    wire N__13301;
    wire N__13300;
    wire N__13299;
    wire N__13296;
    wire N__13295;
    wire N__13294;
    wire N__13293;
    wire N__13292;
    wire N__13285;
    wire N__13282;
    wire N__13275;
    wire N__13270;
    wire N__13267;
    wire N__13262;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13192;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13150;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13108;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13077;
    wire N__13076;
    wire N__13071;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13056;
    wire N__13051;
    wire N__13048;
    wire N__13045;
    wire N__13042;
    wire N__13039;
    wire N__13036;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13006;
    wire N__13005;
    wire N__13004;
    wire N__13001;
    wire N__12996;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12976;
    wire N__12969;
    wire N__12964;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12956;
    wire N__12955;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12937;
    wire N__12936;
    wire N__12935;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12924;
    wire N__12923;
    wire N__12920;
    wire N__12919;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12907;
    wire N__12902;
    wire N__12897;
    wire N__12896;
    wire N__12885;
    wire N__12882;
    wire N__12877;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12816;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12810;
    wire N__12809;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12793;
    wire N__12792;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12772;
    wire N__12769;
    wire N__12766;
    wire N__12763;
    wire N__12758;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12744;
    wire N__12739;
    wire N__12730;
    wire N__12727;
    wire N__12724;
    wire N__12723;
    wire N__12722;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12710;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12690;
    wire N__12689;
    wire N__12688;
    wire N__12687;
    wire N__12686;
    wire N__12685;
    wire N__12680;
    wire N__12679;
    wire N__12674;
    wire N__12671;
    wire N__12670;
    wire N__12667;
    wire N__12666;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12655;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12641;
    wire N__12636;
    wire N__12631;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12615;
    wire N__12610;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12593;
    wire N__12592;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12584;
    wire N__12583;
    wire N__12582;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12567;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12540;
    wire N__12539;
    wire N__12538;
    wire N__12533;
    wire N__12530;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12508;
    wire N__12507;
    wire N__12504;
    wire N__12503;
    wire N__12500;
    wire N__12499;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12448;
    wire N__12447;
    wire N__12442;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12425;
    wire N__12418;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12410;
    wire N__12407;
    wire N__12406;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12343;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12295;
    wire N__12292;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12281;
    wire N__12280;
    wire N__12275;
    wire N__12270;
    wire N__12265;
    wire N__12264;
    wire N__12263;
    wire N__12260;
    wire N__12255;
    wire N__12254;
    wire N__12253;
    wire N__12252;
    wire N__12251;
    wire N__12250;
    wire N__12249;
    wire N__12248;
    wire N__12247;
    wire N__12246;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12217;
    wire N__12216;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12208;
    wire N__12203;
    wire N__12196;
    wire N__12189;
    wire N__12184;
    wire N__12179;
    wire N__12178;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12164;
    wire N__12161;
    wire N__12156;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12034;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12024;
    wire N__12023;
    wire N__12020;
    wire N__12019;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12004;
    wire N__12003;
    wire N__12002;
    wire N__11999;
    wire N__11994;
    wire N__11991;
    wire N__11990;
    wire N__11989;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11966;
    wire N__11963;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11880;
    wire N__11879;
    wire N__11878;
    wire N__11877;
    wire N__11876;
    wire N__11875;
    wire N__11874;
    wire N__11873;
    wire N__11872;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11793;
    wire N__11788;
    wire N__11785;
    wire N__11782;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11770;
    wire N__11767;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11700;
    wire N__11697;
    wire N__11696;
    wire N__11693;
    wire N__11688;
    wire N__11683;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11645;
    wire N__11642;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11623;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11547;
    wire N__11546;
    wire N__11545;
    wire N__11544;
    wire N__11539;
    wire N__11538;
    wire N__11537;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11506;
    wire N__11503;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11457;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11442;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11401;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11389;
    wire N__11386;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11365;
    wire N__11362;
    wire N__11359;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11229;
    wire N__11226;
    wire N__11225;
    wire N__11222;
    wire N__11217;
    wire N__11212;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11193;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11139;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11092;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11058;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11046;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11040;
    wire N__11037;
    wire N__11032;
    wire N__11027;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10985;
    wire N__10978;
    wire N__10977;
    wire N__10976;
    wire N__10975;
    wire N__10974;
    wire N__10971;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10959;
    wire N__10956;
    wire N__10955;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10934;
    wire N__10927;
    wire N__10924;
    wire N__10919;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10894;
    wire N__10891;
    wire N__10890;
    wire N__10887;
    wire N__10884;
    wire N__10883;
    wire N__10882;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10878;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10860;
    wire N__10855;
    wire N__10852;
    wire N__10847;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10831;
    wire N__10828;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10746;
    wire N__10743;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10687;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10664;
    wire N__10663;
    wire N__10662;
    wire N__10659;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10633;
    wire N__10632;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10618;
    wire N__10613;
    wire N__10610;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10584;
    wire N__10575;
    wire N__10568;
    wire N__10563;
    wire N__10552;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10534;
    wire N__10531;
    wire N__10522;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10505;
    wire N__10502;
    wire N__10495;
    wire N__10492;
    wire N__10491;
    wire N__10490;
    wire N__10487;
    wire N__10486;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10468;
    wire N__10465;
    wire N__10456;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10450;
    wire N__10449;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10436;
    wire N__10431;
    wire N__10428;
    wire N__10417;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10411;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10397;
    wire N__10394;
    wire N__10387;
    wire N__10382;
    wire N__10379;
    wire N__10372;
    wire N__10369;
    wire N__10368;
    wire N__10367;
    wire N__10366;
    wire N__10365;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10347;
    wire N__10344;
    wire N__10333;
    wire N__10330;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10322;
    wire N__10321;
    wire N__10316;
    wire N__10313;
    wire N__10312;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10285;
    wire N__10282;
    wire N__10281;
    wire N__10278;
    wire N__10277;
    wire N__10274;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10236;
    wire N__10235;
    wire N__10232;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10188;
    wire N__10183;
    wire N__10180;
    wire N__10179;
    wire N__10176;
    wire N__10175;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10163;
    wire N__10160;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10137;
    wire N__10136;
    wire N__10135;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10120;
    wire N__10111;
    wire N__10110;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10098;
    wire N__10093;
    wire N__10090;
    wire N__10089;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10085;
    wire N__10084;
    wire N__10083;
    wire N__10082;
    wire N__10081;
    wire N__10072;
    wire N__10065;
    wire N__10060;
    wire N__10057;
    wire N__10048;
    wire N__10047;
    wire N__10046;
    wire N__10045;
    wire N__10044;
    wire N__10043;
    wire N__10036;
    wire N__10035;
    wire N__10034;
    wire N__10031;
    wire N__10026;
    wire N__10023;
    wire N__10018;
    wire N__10013;
    wire N__10010;
    wire N__10005;
    wire N__10000;
    wire N__9997;
    wire N__9996;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9933;
    wire N__9932;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9924;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9907;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9882;
    wire N__9877;
    wire N__9862;
    wire N__9859;
    wire N__9858;
    wire N__9857;
    wire N__9856;
    wire N__9855;
    wire N__9852;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9840;
    wire N__9835;
    wire N__9830;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9816;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9808;
    wire N__9805;
    wire N__9804;
    wire N__9803;
    wire N__9800;
    wire N__9789;
    wire N__9784;
    wire N__9783;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9769;
    wire N__9766;
    wire N__9765;
    wire N__9764;
    wire N__9763;
    wire N__9762;
    wire N__9761;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9739;
    wire N__9738;
    wire N__9735;
    wire N__9730;
    wire N__9725;
    wire N__9722;
    wire N__9721;
    wire N__9720;
    wire N__9715;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9699;
    wire N__9698;
    wire N__9695;
    wire N__9690;
    wire N__9685;
    wire N__9682;
    wire N__9677;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9661;
    wire N__9652;
    wire N__9647;
    wire N__9640;
    wire N__9639;
    wire N__9638;
    wire N__9635;
    wire N__9634;
    wire N__9631;
    wire N__9630;
    wire N__9627;
    wire N__9626;
    wire N__9621;
    wire N__9618;
    wire N__9611;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9591;
    wire N__9590;
    wire N__9589;
    wire N__9588;
    wire N__9587;
    wire N__9584;
    wire N__9579;
    wire N__9572;
    wire N__9571;
    wire N__9570;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9551;
    wire N__9546;
    wire N__9545;
    wire N__9544;
    wire N__9543;
    wire N__9542;
    wire N__9541;
    wire N__9540;
    wire N__9539;
    wire N__9538;
    wire N__9537;
    wire N__9536;
    wire N__9535;
    wire N__9530;
    wire N__9521;
    wire N__9512;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9496;
    wire N__9491;
    wire N__9484;
    wire N__9481;
    wire N__9480;
    wire N__9479;
    wire N__9478;
    wire N__9475;
    wire N__9468;
    wire N__9463;
    wire N__9462;
    wire N__9461;
    wire N__9460;
    wire N__9459;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9451;
    wire N__9450;
    wire N__9449;
    wire N__9448;
    wire N__9447;
    wire N__9446;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9427;
    wire N__9422;
    wire N__9413;
    wire N__9408;
    wire N__9405;
    wire N__9404;
    wire N__9403;
    wire N__9400;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9382;
    wire N__9377;
    wire N__9372;
    wire N__9361;
    wire N__9360;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9354;
    wire N__9349;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9337;
    wire N__9334;
    wire N__9325;
    wire N__9324;
    wire N__9323;
    wire N__9322;
    wire N__9319;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9301;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9271;
    wire N__9268;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9240;
    wire N__9237;
    wire N__9226;
    wire N__9223;
    wire N__9222;
    wire N__9221;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9186;
    wire N__9185;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9173;
    wire N__9170;
    wire N__9163;
    wire N__9162;
    wire N__9161;
    wire N__9160;
    wire N__9159;
    wire N__9154;
    wire N__9151;
    wire N__9146;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9024;
    wire N__9023;
    wire N__9022;
    wire N__9021;
    wire N__9016;
    wire N__9013;
    wire N__9008;
    wire N__9001;
    wire N__9000;
    wire N__8995;
    wire N__8992;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8970;
    wire N__8969;
    wire N__8968;
    wire N__8967;
    wire N__8966;
    wire N__8959;
    wire N__8952;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8940;
    wire N__8939;
    wire N__8938;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8923;
    wire N__8918;
    wire N__8911;
    wire N__8910;
    wire N__8909;
    wire N__8908;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8895;
    wire N__8894;
    wire N__8893;
    wire N__8890;
    wire N__8883;
    wire N__8880;
    wire N__8869;
    wire N__8860;
    wire N__8859;
    wire N__8858;
    wire N__8855;
    wire N__8854;
    wire N__8853;
    wire N__8852;
    wire N__8851;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8839;
    wire N__8836;
    wire N__8829;
    wire N__8818;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8806;
    wire N__8803;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8748;
    wire N__8745;
    wire N__8740;
    wire N__8737;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8701;
    wire N__8700;
    wire N__8699;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8671;
    wire N__8668;
    wire N__8665;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8646;
    wire N__8645;
    wire N__8644;
    wire N__8643;
    wire N__8642;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8630;
    wire N__8629;
    wire N__8626;
    wire N__8621;
    wire N__8620;
    wire N__8617;
    wire N__8612;
    wire N__8609;
    wire N__8608;
    wire N__8607;
    wire N__8602;
    wire N__8601;
    wire N__8600;
    wire N__8599;
    wire N__8596;
    wire N__8589;
    wire N__8584;
    wire N__8581;
    wire N__8574;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8547;
    wire N__8546;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8523;
    wire N__8522;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8506;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8488;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8478;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8457;
    wire N__8456;
    wire N__8455;
    wire N__8446;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8433;
    wire N__8428;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8410;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8367;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8350;
    wire N__8349;
    wire N__8348;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8323;
    wire N__8320;
    wire N__8319;
    wire N__8318;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8265;
    wire N__8264;
    wire N__8263;
    wire N__8258;
    wire N__8253;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8227;
    wire N__8224;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8203;
    wire N__8202;
    wire N__8201;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8185;
    wire N__8184;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8157;
    wire N__8154;
    wire N__8153;
    wire N__8152;
    wire N__8149;
    wire N__8144;
    wire N__8141;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8124;
    wire N__8121;
    wire N__8118;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8079;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8064;
    wire N__8063;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8049;
    wire N__8048;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7978;
    wire N__7977;
    wire N__7976;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7964;
    wire N__7961;
    wire N__7956;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7939;
    wire N__7938;
    wire N__7937;
    wire N__7936;
    wire N__7933;
    wire N__7926;
    wire N__7925;
    wire N__7924;
    wire N__7923;
    wire N__7922;
    wire N__7917;
    wire N__7912;
    wire N__7911;
    wire N__7910;
    wire N__7907;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7887;
    wire N__7876;
    wire N__7875;
    wire N__7874;
    wire N__7873;
    wire N__7872;
    wire N__7871;
    wire N__7870;
    wire N__7867;
    wire N__7860;
    wire N__7853;
    wire N__7852;
    wire N__7845;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7828;
    wire N__7825;
    wire N__7824;
    wire N__7823;
    wire N__7820;
    wire N__7819;
    wire N__7818;
    wire N__7817;
    wire N__7816;
    wire N__7811;
    wire N__7810;
    wire N__7809;
    wire N__7806;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7747;
    wire N__7744;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7710;
    wire N__7709;
    wire N__7708;
    wire N__7705;
    wire N__7702;
    wire N__7697;
    wire N__7690;
    wire N__7689;
    wire N__7684;
    wire N__7683;
    wire N__7682;
    wire N__7681;
    wire N__7678;
    wire N__7673;
    wire N__7670;
    wire N__7665;
    wire N__7664;
    wire N__7663;
    wire N__7662;
    wire N__7659;
    wire N__7656;
    wire N__7651;
    wire N__7648;
    wire N__7639;
    wire N__7638;
    wire N__7635;
    wire N__7634;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7619;
    wire N__7612;
    wire N__7609;
    wire N__7608;
    wire N__7607;
    wire N__7606;
    wire N__7601;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7590;
    wire N__7589;
    wire N__7588;
    wire N__7585;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7569;
    wire N__7558;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7539;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7516;
    wire N__7513;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7485;
    wire N__7484;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7472;
    wire N__7469;
    wire N__7462;
    wire N__7461;
    wire N__7456;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7437;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7395;
    wire N__7392;
    wire N__7391;
    wire N__7388;
    wire N__7387;
    wire N__7386;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7366;
    wire N__7363;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7347;
    wire N__7346;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7332;
    wire N__7331;
    wire N__7326;
    wire N__7323;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7293;
    wire N__7290;
    wire N__7289;
    wire N__7288;
    wire N__7287;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7267;
    wire N__7264;
    wire N__7261;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7204;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7192;
    wire N__7191;
    wire N__7188;
    wire N__7183;
    wire N__7180;
    wire N__7177;
    wire N__7174;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7162;
    wire N__7159;
    wire N__7156;
    wire N__7153;
    wire N__7150;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7107;
    wire N__7106;
    wire N__7103;
    wire N__7102;
    wire N__7101;
    wire N__7098;
    wire N__7089;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7077;
    wire N__7074;
    wire N__7071;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7008;
    wire N__7007;
    wire N__7004;
    wire N__7003;
    wire N__7000;
    wire N__6999;
    wire N__6996;
    wire N__6987;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6942;
    wire N__6939;
    wire N__6938;
    wire N__6937;
    wire N__6930;
    wire N__6927;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6796;
    wire N__6793;
    wire N__6790;
    wire N__6787;
    wire N__6784;
    wire N__6781;
    wire \Clock50MHz.PixelClock ;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_6_0_;
    wire un21_beamy_cry_1;
    wire un21_beamy_cry_2;
    wire un21_beamy_cry_3;
    wire un21_beamy_cry_4;
    wire un21_beamy_cry_5;
    wire un21_beamy_cry_6;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire bfn_1_7_0_;
    wire bfn_1_8_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOGZ0Z53;
    wire bfn_1_9_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOSZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRSZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LKZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01_cascade_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0;
    wire bfn_1_10_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOLZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IGZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMGZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0;
    wire bfn_1_11_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICMZ0Z321;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPMZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KHZ0Z2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0;
    wire bfn_1_12_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CRZ0Z2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGIZ0Z3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJZ0Z6874;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7;
    wire un21_beamy_cry_4_c_RNIGUAZ0Z3;
    wire un21_beamy_cry_6_c_RNIK4DZ0Z3;
    wire beamY_fastZ0Z_7;
    wire beamY_fastZ0Z_5;
    wire un21_beamy_cry_1_c_RNIALZ0Z73;
    wire un5_visibley_c6_0_0_0;
    wire beamY_fast_RNI35GAZ0Z_2_cascade_;
    wire un21_beamy_cry_2_c_RNICOZ0Z83;
    wire bfn_2_7_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2;
    wire bfn_2_8_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2LZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RCZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5;
    wire beamY_RNIFJ0L_0Z0Z_8;
    wire beamY_RNI19IJ_0Z0Z_9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7;
    wire beamY_i_2_cascade_;
    wire un114_pixel_1_0_3__chessboardpixel_un200_pixellto4Z0Z_1_cascade_;
    wire chessboardpixel_un200_pixellt10_cascade_;
    wire chessboardpixel_un200_pixel_0_1_cascade_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5;
    wire beamY_i_2;
    wire bfn_2_10_0_;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81BZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEGZ0Z5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODGZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87VZ0Z68;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4JZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05UZ0Z8;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGKZ0;
    wire chessboardpixel_un174_pixel_0_1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0;
    wire bfn_2_11_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHFZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJZ0Z5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0;
    wire un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1Z0Z_1;
    wire un114_pixel_1_0_3__un1_beamylto9Z0Z_0_cascade_;
    wire un4_beamylt6_cascade_;
    wire un5_visibley_ac0_11_d;
    wire un5_visibley_ac0_11_0_1;
    wire un114_pixel_1_0_3__un1_beamylto9_3;
    wire beamY_fastZ0Z_2;
    wire beamYZ0Z_5;
    wire beamY_fastZ0Z_3;
    wire beamY_fast_RNIM4P7Z0Z_2_cascade_;
    wire beamYZ0Z_6;
    wire un5_visibley_c5;
    wire un5_visibley_c5_cascade_;
    wire un114_pixel_1_0_3__un5_beamxZ0Z_5_cascade_;
    wire un114_pixel_1_0_3__g0_1Z0Z_0_cascade_;
    wire un4_beamylt8_0;
    wire un5_visibley_c2;
    wire un1_beamy_4;
    wire beamYZ0Z_8;
    wire beamYZ0Z_9;
    wire un114_pixel_1_0_3__un8_beamylto9Z0Z_1_cascade_;
    wire beamYZ0Z_7;
    wire row_1_if_generate_plus_mult1_un75_sum_cZ0Z4;
    wire row_1_if_generate_plus_mult1_un75_sum_cZ0Z4_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_;
    wire row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1;
    wire row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_;
    wire if_generate_plus_mult1_un68_sum_axbxc3;
    wire row_1_if_generate_plus_mult1_un68_sum_c5_0_nsZ0Z_1;
    wire row_1_if_generate_plus_mult1_un68_sum_c5;
    wire row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5;
    wire if_generate_plus_mult1_un54_sum_axbxc3;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_c5;
    wire row_1_if_generate_plus_mult1_un61_sum_c5_cascade_;
    wire row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0;
    wire if_generate_plus_mult1_un68_sum_c5_0_bm;
    wire row_1_if_generate_plus_mult1_un61_sum_ac0_7_c;
    wire bfn_4_11_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KCZ0Z4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGSZ0Z6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8;
    wire bfn_4_13_0_;
    wire counter_cry_1;
    wire counter_cry_2;
    wire counter_cry_3;
    wire counter_cry_4;
    wire slaveselect_1_0_4_cascade_;
    wire counter_30;
    wire un3_slaveselect_cascade_;
    wire counter_29;
    wire counter_31_cascade_;
    wire counterZ0Z_0;
    wire counterZ0Z_3;
    wire counterZ0Z_1;
    wire un1_counterlto3_0_cascade_;
    wire counterZ0Z_2;
    wire g0_0_1_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_c5;
    wire un5_visibley_0_29;
    wire chary_if_generate_plus_mult1_un61_sum_c5_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_0_1_5;
    wire chary_if_generate_plus_mult1_un68_sum_c4_0_cascade_;
    wire g0_0_3;
    wire g1_0_cascade_;
    wire un4_beamylt6;
    wire chary_if_generate_plus_mult1_un75_sum_c5_N_9_cascade_;
    wire g0_1_2;
    wire g0_2_0;
    wire chary_if_generate_plus_mult1_un61_sum_1_0_1_0_3;
    wire beamY_RNINITP61Z0Z_5_cascade_;
    wire beamY_RNINITP61_1Z0Z_5;
    wire chary_if_generate_plus_mult1_un40_sum_axb3;
    wire chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0_cascade_;
    wire chary_if_generate_plus_mult1_un47_sum_axbxc5_2;
    wire chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_;
    wire chary_if_generate_plus_mult1_un40_sum_c4;
    wire chary_if_generate_plus_mult1_un47_sum_c5;
    wire beamY_RNITURI3_0Z0Z_7_cascade_;
    wire beamY_RNITURI3Z0Z_7;
    wire un4_beamy_0;
    wire un8_beamy;
    wire un114_pixel_1_0_3__un15_beamyZ0Z_2;
    wire un1_beamx_2_cascade_;
    wire un114_pixel_1_0_3__un5_beamxZ0Z_3;
    wire beamYZ0Z_4;
    wire un114_pixel_1_0_3__g0_1Z0Z_3;
    wire un114_pixel_1_0_3__un18_beamylto9Z0Z_2_cascade_;
    wire un18_beamylt10_0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum;
    wire un13_beamylt7;
    wire if_generate_plus_mult1_un75_sum_axbxc5;
    wire if_generate_plus_mult1_un75_sum_axbxc3;
    wire row_1_if_generate_plus_mult1_un82_sum_axb4_i_cascade_;
    wire row_1_if_generate_plus_mult1_un82_sum_ac0_7_0Z0Z_1;
    wire bfn_5_9_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_5_10_0_;
    wire un8_beamx_cry_9;
    wire row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0;
    wire bfn_5_11_0_;
    wire charx_if_generate_plus_mult1_un19_sum_cry_2;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i;
    wire counter_27;
    wire counterZ0Z_5;
    wire slaveselect_1_0_4;
    wire un1_slaveselect_1_i;
    wire un3_slaveselect;
    wire counter_28;
    wire counterZ0Z_4;
    wire slaveselectZ0;
    wire un1_counter_0;
    wire nCS1_c;
    wire nCS1_0_sqmuxa;
    wire beamY_RNI2TEJF4Z0Z_4_cascade_;
    wire un114_pixel_1_0_3__g0_8Z0Z_1;
    wire chary_if_generate_plus_mult1_un61_sum_0_3_cascade_;
    wire un114_pixel_1_0_3__g0_1Z0Z_1_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_0_3;
    wire un114_pixel_1_0_3__g0_3Z0Z_0_cascade_;
    wire chary_if_generate_plus_mult1_un75_sum_i_0_5;
    wire chary_if_generate_plus_mult1_un68_sum_c4_0;
    wire un114_pixel_1_0_3__g0Z0Z_1_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_0_0_0_0_5;
    wire g2;
    wire un114_pixel_1_0_3__g0Z0Z_3_cascade_;
    wire beamY_RNITFRN03Z0Z_5;
    wire chary_if_generate_plus_mult1_un75_sum_c5;
    wire beamY_RNIH9THADZ0Z_4_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_axb3_0;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_d;
    wire beamY_RNIKHPCA1Z0Z_4;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_d_cascade_;
    wire chary_if_generate_plus_mult1_un68_sum_axb4;
    wire beamY_RNI2TEJF4Z0Z_4;
    wire chary_if_generate_plus_mult1_un68_sum_c4;
    wire chary_if_generate_plus_mult1_un61_sum_axb4_0;
    wire g0_0_x2_1_1_cascade_;
    wire g0_3_2;
    wire beamY_RNIARUFBZ0Z_5_cascade_;
    wire beamY_RNIGS0LBZ0Z_5;
    wire chary_if_generate_plus_mult1_un54_sum_c5;
    wire chary_if_generate_plus_mult1_un54_sum_c5_cascade_;
    wire chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0;
    wire chary_if_generate_plus_mult1_un61_sum_axb3_0_0;
    wire beamY_RNIDO3IZ0Z_9;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum;
    wire chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0;
    wire g0_4_2;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum;
    wire chary_if_generate_plus_mult1_un54_sum_axb3;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum;
    wire chary_if_generate_plus_mult1_un54_sum_axbxc5_1;
    wire beamY_RNI2MTA1Z0Z_9;
    wire chary_if_generate_plus_mult1_un54_sum_c4_cascade_;
    wire beamY_RNICG8P9Z0Z_7;
    wire chary_if_generate_plus_mult1_un61_sum_axbxc5_1;
    wire un3_beamx_0_cascade_;
    wire un1_beamx_2;
    wire HSync_c;
    wire bfn_6_8_0_;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2;
    wire charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8VZ0;
    wire charx_if_generate_plus_mult1_un26_sum_cry_3;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4;
    wire un1_beamxlt10_0;
    wire beamXZ0Z_10;
    wire un114_pixel_1_0_3__un3_beamxZ0Z_5_cascade_;
    wire un114_pixel_1_0_3__un3_beamxZ0Z_7;
    wire un18_beamylt4;
    wire charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO;
    wire charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKFZ0;
    wire charx_if_generate_plus_mult1_un19_sum_i;
    wire bfn_6_10_0_;
    wire beamXZ0Z_1;
    wire un5_visiblex_cry_0;
    wire beamXZ0Z_2;
    wire un5_visiblex_cry_1;
    wire beamXZ0Z_3;
    wire un5_visiblex_cry_2;
    wire beamXZ0Z_4;
    wire un5_visiblex_cry_3;
    wire beamXZ0Z_5;
    wire un5_visiblex_cry_4;
    wire beamXZ0Z_6;
    wire un5_visiblex_cry_5;
    wire beamXZ0Z_7;
    wire un5_visiblex_cry_6;
    wire un5_visiblex_cry_7;
    wire beamXZ0Z_8;
    wire bfn_6_11_0_;
    wire beamXZ0Z_9;
    wire un5_visiblex_cry_8;
    wire un116_pixel_3_bm_2_cascade_;
    wire un114_pixel_1_0_3__N_5_1_0;
    wire un114_pixel_1_0_3__un116_pixel_4_ns_1_0_7_cascade_;
    wire un114_pixel_1_0_3__g2_1Z0Z_0;
    wire beamY_RNIH9THADZ0Z_4;
    wire beamYZ0Z_3;
    wire N_345_0_0_1;
    wire font_un28_pixel_29_cascade_;
    wire un116_pixel_5_am_6_cascade_;
    wire g1_1;
    wire g0_0_x2_1;
    wire un114_pixel_1_0_3__un116_pixel_2_ns_1Z0Z_2_cascade_;
    wire un114_pixel_1_0_3__un116_pixel_5_ns_1Z0Z_2_cascade_;
    wire un116_pixel_5_ns_1Z0Z_4_cascade_;
    wire un116_pixel_5_ns_2;
    wire N_362;
    wire un116_pixel_7_ns_1_6_cascade_;
    wire N_379;
    wire un116_pixel_3_ns_2;
    wire beamY_RNI57H3N31_0Z0Z_1_cascade_;
    wire beamY_RNI896FQ3Z0Z_0;
    wire beamY_RNI896FQ3Z0Z_0_cascade_;
    wire beamY_RNI57H3N31Z0Z_1;
    wire un116_pixel_2_ns_1_0_6_cascade_;
    wire beamY_RNIGO5PPVZ0Z_0;
    wire N_41;
    wire un3_beamx_0;
    wire un5_beamx_0;
    wire bfn_7_7_0_;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_1;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un68_sum_cry_4;
    wire column_1_if_generate_plus_mult1_un61_sum_iZ0;
    wire row_1_if_generate_plus_mult1_un54_sum_cZ0Z5;
    wire un5_rowlto3_i;
    wire bfn_7_8_0_;
    wire N_575_i;
    wire if_generate_plus_mult1_un61_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_1;
    wire if_generate_plus_mult1_un61_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un61_sum_cry_4;
    wire column_1_if_generate_plus_mult1_un54_sum_i_5;
    wire bfn_7_9_0_;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1;
    wire charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2;
    wire charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HLZ0;
    wire charx_if_generate_plus_mult1_un33_sum_cry_3;
    wire charx_if_generate_plus_mult1_un33_sum_axb_5;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4;
    wire charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5;
    wire charx_if_generate_plus_mult1_un26_sum_i_5;
    wire bfn_7_10_0_;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1;
    wire charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072;
    wire charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2;
    wire charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0;
    wire charx_if_generate_plus_mult1_un33_sum_i_5;
    wire charx_if_generate_plus_mult1_un40_sum_cry_3;
    wire charx_if_generate_plus_mult1_un40_sum_axb_5;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4;
    wire charx_if_generate_plus_mult1_un33_sum_i;
    wire charx_if_generate_plus_mult1_un26_sum_i;
    wire bfn_7_11_0_;
    wire if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_1;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_2;
    wire N_204_0_i;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_3;
    wire column_1_if_generate_plus_mult1_un47_sum_0_cry_4;
    wire un5_visiblex_i_25;
    wire if_generate_plus_mult1_un47_sum_0_cry_3_ma;
    wire if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx;
    wire bfn_7_12_0_;
    wire if_generate_plus_mult1_un54_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_1;
    wire if_generate_plus_mult1_un54_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un54_sum_cry_4;
    wire column_1_if_generate_plus_mult1_un47_sum0_3;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_;
    wire if_generate_plus_mult1_un54_sum_axb_4_l_fx;
    wire bfn_7_13_0_;
    wire charx_if_generate_plus_mult1_un40_sum_i;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1;
    wire charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3;
    wire charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEBZ0Z2;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2;
    wire charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLITZ0Z2;
    wire charx_if_generate_plus_mult1_un40_sum_i_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_3;
    wire charx_if_generate_plus_mult1_un47_sum_axb_5;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6_cascade_;
    wire charx_if_generate_plus_mult1_un47_sum;
    wire bfn_7_14_0_;
    wire charx_if_generate_plus_mult1_un47_sum_i;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1;
    wire charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6;
    wire charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0OZ0Z3;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2;
    wire charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCDZ0Z16;
    wire charx_if_generate_plus_mult1_un47_sum_i_5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_3;
    wire charx_if_generate_plus_mult1_un54_sum_axb_5;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4;
    wire charx_if_generate_plus_mult1_un54_sum;
    wire bfn_7_15_0_;
    wire charx_if_generate_plus_mult1_un54_sum_i;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1;
    wire charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLMZ0Z67;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2;
    wire charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSAZ0;
    wire charx_if_generate_plus_mult1_un61_sum_cry_3;
    wire charx_if_generate_plus_mult1_un61_sum_axb_5;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0_cascade_;
    wire charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0;
    wire charx_if_generate_plus_mult1_un54_sum_i_5;
    wire VSync_c;
    wire un116_pixel_3_am_2;
    wire N_1556_0_cascade_;
    wire N_347_0;
    wire font_un28_pixel_0_29;
    wire N_368_0;
    wire un114_pixel_1_0_3__font_un126_pixel_1_d_ns_1_0_cascade_;
    wire N_389_0;
    wire N_346_0_0_1;
    wire g0_cascade_;
    wire N_36_cascade_;
    wire un116_pixel_3_ns_1_1_cascade_;
    wire font_un3_pixel_29_cascade_;
    wire un116_pixel_5_bm_6;
    wire un116_pixel_4_bm_1;
    wire beamY_RNI1C50FS3Z0Z_0_cascade_;
    wire un116_pixel_3_bm_1_6_cascade_;
    wire beamY_RNIOHI2NGZ0Z_0;
    wire N_364_cascade_;
    wire un116_pixel_7_ns_1_4_cascade_;
    wire beamY_RNI2L0T663Z0Z_0;
    wire column_0111_1_0;
    wire beamY_RNI1J75181Z0Z_1;
    wire font_un126_pixel_6_am_cascade_;
    wire un1_beamy_0;
    wire N_1075_0_cascade_;
    wire N_400;
    wire Pixel_r_rn_0_cascade_;
    wire Pixel_c;
    wire PixelClock_g;
    wire font_un28_pixel_0_0_29;
    wire font_un126_pixel_2_bm;
    wire un114_pixel_1_0_3__font_un126_pixel_7_d_ns_1_0_0;
    wire beamY_RNIHHB5F01Z0Z_4;
    wire beamYZ0Z_2;
    wire beamY_RNI7OE17CZ0Z_0;
    wire beamY_RNIVU1O9RZ0Z_1;
    wire font_un126_pixel_6_bm;
    wire charx_if_generate_plus_mult1_un1_sum_axb1_cascade_;
    wire un15_beamy;
    wire r_i1_mux_cascade_;
    wire un114_pixel_1_0_3__font_un126_pixel_mZ0Z_1_cascade_;
    wire chary_24;
    wire un114_pixel_1_0_3__font_un126_pixel_m_1_0_cascade_;
    wire chary_23;
    wire un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3;
    wire un1_beamylto9;
    wire un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3_cascade_;
    wire Pixel_r_sn;
    wire beamXZ0Z_0;
    wire un114_pixel_1_0_3__font_un57_pixelZ0Z_0;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum;
    wire if_generate_plus_mult1_un61_sum_axbxc5;
    wire un114_pixel_1_0_3__un4_row_8Z0Z_3_cascade_;
    wire un114_pixel_1_0_3__un4_row_8_7Z0Z_1;
    wire chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum;
    wire chary_if_generate_plus_mult1_un33_sum_axb3;
    wire if_generate_plus_mult1_un54_sum_s_5;
    wire un114_pixel_1_0_3__un4_row_8Z0Z_2;
    wire row_1_if_generate_plus_mult1_un75_sum_cZ0Z5;
    wire if_generate_plus_mult1_un68_sum_axbxc5;
    wire row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2;
    wire un114_pixel_1_0_3__un4_row_8Z0Z_7;
    wire un114_pixel_1_0_3__un4_rowZ0Z_8;
    wire row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1;
    wire row_1_if_generate_plus_mult1_un82_sum_c5;
    wire un114_pixel_1_0_3__un4_rowZ0Z_8_cascade_;
    wire un114_pixel_1_0_3__Pixel_3_sqmuxaZ0Z_0;
    wire Pixel_3_sqmuxa;
    wire bfn_8_10_0_;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4_c_invZ0;
    wire charx_if_generate_plus_mult1_un75_sum_cry_3;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843_cascade_;
    wire charx_if_generate_plus_mult1_un68_sum_i;
    wire un114_pixel_1_0_3__un4_row_8Z0Z_0;
    wire charx_if_generate_plus_mult1_un68_sum_i_5;
    wire if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx;
    wire column_1_if_generate_plus_mult1_un54_sum_axb_2_sxZ0_cascade_;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2_cascade_;
    wire if_generate_plus_mult1_un54_sum_axb_2_l_fx;
    wire column_1_if_generate_plus_mult1_un47_sum0_4;
    wire if_generate_plus_mult1_un47_sum_m_5_cascade_;
    wire column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un47_sum0_2;
    wire if_generate_plus_mult1_un47_sum_m_5;
    wire if_generate_plus_mult1_un54_sum_axb_3_l_fx;
    wire column_1_if_generate_plus_mult1_un47_sum0_5;
    wire N_584_i;
    wire N_37_i;
    wire bfn_8_14_0_;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5RZ0;
    wire charx_if_generate_plus_mult1_un68_sum_cry_1;
    wire charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0;
    wire charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRDZ0;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BVZ0Z81;
    wire charx_if_generate_plus_mult1_un68_sum_cry_2;
    wire charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0LZ0;
    wire charx_if_generate_plus_mult1_un61_sum_i_5;
    wire charx_if_generate_plus_mult1_un75_sum_axb_5;
    wire charx_if_generate_plus_mult1_un68_sum_cry_3;
    wire charx_if_generate_plus_mult1_un68_sum_axb_5;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4;
    wire charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1;
    wire charx_if_generate_plus_mult1_un61_sum_i;
    wire N_41_0;
    wire column_0111_0;
    wire un116_pixel_3_ns_1_0_3;
    wire un114_pixel_1_0_3__g1Z0Z_4;
    wire N_1583_0_cascade_;
    wire N_26_0_0;
    wire un116_pixel_2_amZ0Z_1_cascade_;
    wire un116_pixel_6_1;
    wire column_0001_0_cascade_;
    wire beamY_RNILBST4T2Z0Z_1;
    wire beamY_RNIT81CMJ2Z0Z_1_cascade_;
    wire font_un126_pixel_2_am;
    wire un116_pixel_4_am_1;
    wire N_36;
    wire un116_pixel_5_amZ0Z_5;
    wire un116_pixel_2_amZ0Z_5;
    wire N_385;
    wire N_325;
    wire un116_pixel_2_bmZ0Z_1;
    wire un114_pixel_1_0_3__un116_pixel_6_1Z0Z_1;
    wire un116_pixel_1_4;
    wire N_374_0;
    wire font_un3_pixel_29;
    wire un116_pixel_7_x0_0_cascade_;
    wire un116_pixel_7_x1_0;
    wire un116_pixel_7_ns_0;
    wire un116_pixel_2_bm_0;
    wire un114_pixel_1_0_3__un116_pixel_5_ns_1_0Z0Z_0;
    wire chessboardpixel_un152_pixel_24;
    wire un114_pixel_1_0_3__un116_pixel_6_1_1Z0Z_1;
    wire charx_if_generate_plus_mult1_un1_sum_axb1;
    wire bfn_9_8_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3EZ0Z987;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0;
    wire bfn_9_9_0_;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8TZ0Z77;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1;
    wire font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4;
    wire font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77Z0Z_0;
    wire charx_i_23;
    wire charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1;
    wire charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2;
    wire charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843;
    wire charx_i_24;
    wire bfn_9_11_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUHZ0Z2;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIVZ0Z6153;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i;
    wire charx_if_generate_plus_mult1_un40_sum;
    wire bfn_9_12_0_;
    wire un5_visiblex_i_0_25;
    wire column_1_if_generate_plus_mult1_un47_sum1_2;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_1;
    wire if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx;
    wire N_858_i;
    wire column_1_if_generate_plus_mult1_un47_sum1_3;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_2;
    wire if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx;
    wire column_1_if_generate_plus_mult1_un47_sum1_4;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_3;
    wire column_1_if_generate_plus_mult1_un47_sum_1_cry_4;
    wire column_1_if_generate_plus_mult1_un47_sum1_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8;
    wire charx_if_generate_plus_mult1_un33_sum;
    wire N_66;
    wire bfn_9_13_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5LZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7JZ0Z31;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i;
    wire Clock12MHz_c_g;
    wire GB_BUFFER_Clock12MHz_c_g_THRU_CO;
    wire N_1557_0;
    wire N_41_0_0_0;
    wire N_563;
    wire un116_pixel_5_bmZ0Z_5_cascade_;
    wire un116_pixel_6_ns_1_5;
    wire un116_pixel_2_bmZ0Z_5;
    wire un114_pixel_7_1_7__N_9_cascade_;
    wire un114_pixel_1_0_3__un116_pixel_3_ns_1Z0Z_0_cascade_;
    wire un114_pixel_6_1_5__N_8;
    wire N_371;
    wire beamY_RNIJUCG3J3Z0Z_1;
    wire charx_if_generate_plus_mult1_un75_sum;
    wire bfn_11_6_0_;
    wire G_345;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_1;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_2;
    wire G_346;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un82_sum_cry_4;
    wire un5_rowlto0_cascade_;
    wire un116_pixel_1_bmZ0Z_1;
    wire beamYZ0Z_1;
    wire un116_pixel_1_bmZ0Z_1_cascade_;
    wire beamY_RNIV622TRZ0Z_1;
    wire un116_pixel_2_ns_1_4;
    wire beamYZ0Z_0;
    wire beamY_RNIITCG3J3Z0Z_0;
    wire bfn_11_7_0_;
    wire column_1_if_generate_plus_mult1_un68_sum_iZ0;
    wire if_generate_plus_mult1_un75_sum_cry_2_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_1;
    wire if_generate_plus_mult1_un68_sum_cry_2_s;
    wire if_generate_plus_mult1_un75_sum_cry_3_s;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_2;
    wire column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_3;
    wire column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5;
    wire column_1_if_generate_plus_mult1_un75_sum_cry_4;
    wire un5_rowlto1;
    wire un5_rowlto0;
    wire un5_rowlto1_cascade_;
    wire un5_rowlto3;
    wire un116_pixel_2_am_0;
    wire if_generate_plus_mult1_un68_sum_cry_3_s;
    wire if_generate_plus_mult1_un75_sum_axb_4_l_fx;
    wire un5_rowlto2;
    wire un5_rowlto2_i;
    wire charx_if_generate_plus_mult1_un68_sum;
    wire column_1_if_generate_plus_mult1_un75_sum_iZ0;
    wire bfn_11_11_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire charx_if_generate_plus_mult1_un26_sum;
    wire bfn_11_12_0_;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHGZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire CONSTANT_ONE_NET;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6QZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0;
    wire CO3_0;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKNZ0;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__14306),
            .RESETB(N__16348),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    PRE_IO_GBUF Clock12MHz_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__16511),
            .GLOBALBUFFEROUTPUT(Clock12MHz_c_g));
    defparam Clock12MHz_ibuf_gb_io_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_gb_io_iopad (
            .OE(N__16513),
            .DIN(N__16512),
            .DOUT(N__16511),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_gb_io_preio (
            .PADOEN(N__16513),
            .PADOUT(N__16512),
            .PADIN(N__16511),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__16502),
            .DIN(N__16501),
            .DOUT(N__16500),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__16502),
            .PADOUT(N__16501),
            .PADIN(N__16500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11668),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__16493),
            .DIN(N__16492),
            .DOUT(N__16491),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__16493),
            .PADOUT(N__16492),
            .PADIN(N__16491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam nCS1_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD nCS1_obuf_iopad (
            .OE(N__16484),
            .DIN(N__16483),
            .DOUT(N__16482),
            .PACKAGEPIN(nCS1));
    defparam nCS1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCS1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCS1_obuf_preio (
            .PADOEN(N__16484),
            .PADOUT(N__16483),
            .PADIN(N__16482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8818),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__16475),
            .DIN(N__16474),
            .DOUT(N__16473),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__16475),
            .PADOUT(N__16474),
            .PADIN(N__16473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11896),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam nCS2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD nCS2_obuf_iopad (
            .OE(N__16466),
            .DIN(N__16465),
            .DOUT(N__16464),
            .PACKAGEPIN(nCS2));
    defparam nCS2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam nCS2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO nCS2_obuf_preio (
            .PADOEN(N__16466),
            .PADOUT(N__16465),
            .PADIN(N__16464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8817),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SCLK1_obuft_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SCLK1_obuft_iopad (
            .OE(N__16457),
            .DIN(N__16456),
            .DOUT(N__16455),
            .PACKAGEPIN(SCLK1));
    defparam SCLK1_obuft_preio.NEG_TRIGGER=1'b0;
    defparam SCLK1_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO SCLK1_obuft_preio (
            .PADOEN(N__16457),
            .PADOUT(N__16456),
            .PADIN(N__16455),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8992),
            .DIN0(),
            .DOUT0(N__14308),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam SCLK2_obuft_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD SCLK2_obuft_iopad (
            .OE(N__16448),
            .DIN(N__16447),
            .DOUT(N__16446),
            .PACKAGEPIN(SCLK2));
    defparam SCLK2_obuft_preio.NEG_TRIGGER=1'b0;
    defparam SCLK2_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO SCLK2_obuft_preio (
            .PADOEN(N__16448),
            .PADOUT(N__16447),
            .PADIN(N__16446),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8991),
            .DIN0(),
            .DOUT0(N__14307),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__3800 (
            .O(N__16429),
            .I(N__16426));
    InMux I__3799 (
            .O(N__16426),
            .I(N__16423));
    LocalMux I__3798 (
            .O(N__16423),
            .I(N__16420));
    Span4Mux_h I__3797 (
            .O(N__16420),
            .I(N__16417));
    Odrv4 I__3796 (
            .O(N__16417),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHGZ0));
    InMux I__3795 (
            .O(N__16414),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__3794 (
            .O(N__16411),
            .I(N__16408));
    InMux I__3793 (
            .O(N__16408),
            .I(N__16404));
    CascadeMux I__3792 (
            .O(N__16407),
            .I(N__16398));
    LocalMux I__3791 (
            .O(N__16404),
            .I(N__16391));
    CascadeMux I__3790 (
            .O(N__16403),
            .I(N__16388));
    CascadeMux I__3789 (
            .O(N__16402),
            .I(N__16385));
    InMux I__3788 (
            .O(N__16401),
            .I(N__16380));
    InMux I__3787 (
            .O(N__16398),
            .I(N__16377));
    InMux I__3786 (
            .O(N__16397),
            .I(N__16374));
    InMux I__3785 (
            .O(N__16396),
            .I(N__16371));
    InMux I__3784 (
            .O(N__16395),
            .I(N__16368));
    InMux I__3783 (
            .O(N__16394),
            .I(N__16365));
    Span4Mux_v I__3782 (
            .O(N__16391),
            .I(N__16361));
    InMux I__3781 (
            .O(N__16388),
            .I(N__16356));
    InMux I__3780 (
            .O(N__16385),
            .I(N__16356));
    CascadeMux I__3779 (
            .O(N__16384),
            .I(N__16352));
    CascadeMux I__3778 (
            .O(N__16383),
            .I(N__16349));
    LocalMux I__3777 (
            .O(N__16380),
            .I(N__16343));
    LocalMux I__3776 (
            .O(N__16377),
            .I(N__16343));
    LocalMux I__3775 (
            .O(N__16374),
            .I(N__16340));
    LocalMux I__3774 (
            .O(N__16371),
            .I(N__16333));
    LocalMux I__3773 (
            .O(N__16368),
            .I(N__16333));
    LocalMux I__3772 (
            .O(N__16365),
            .I(N__16333));
    InMux I__3771 (
            .O(N__16364),
            .I(N__16330));
    Sp12to4 I__3770 (
            .O(N__16361),
            .I(N__16327));
    LocalMux I__3769 (
            .O(N__16356),
            .I(N__16324));
    InMux I__3768 (
            .O(N__16355),
            .I(N__16319));
    InMux I__3767 (
            .O(N__16352),
            .I(N__16319));
    InMux I__3766 (
            .O(N__16349),
            .I(N__16316));
    IoInMux I__3765 (
            .O(N__16348),
            .I(N__16313));
    Span4Mux_v I__3764 (
            .O(N__16343),
            .I(N__16310));
    Span4Mux_h I__3763 (
            .O(N__16340),
            .I(N__16303));
    Span4Mux_v I__3762 (
            .O(N__16333),
            .I(N__16303));
    LocalMux I__3761 (
            .O(N__16330),
            .I(N__16303));
    Span12Mux_s10_h I__3760 (
            .O(N__16327),
            .I(N__16294));
    Sp12to4 I__3759 (
            .O(N__16324),
            .I(N__16294));
    LocalMux I__3758 (
            .O(N__16319),
            .I(N__16294));
    LocalMux I__3757 (
            .O(N__16316),
            .I(N__16294));
    LocalMux I__3756 (
            .O(N__16313),
            .I(N__16291));
    Span4Mux_h I__3755 (
            .O(N__16310),
            .I(N__16286));
    Span4Mux_v I__3754 (
            .O(N__16303),
            .I(N__16286));
    Span12Mux_v I__3753 (
            .O(N__16294),
            .I(N__16281));
    Span12Mux_s1_v I__3752 (
            .O(N__16291),
            .I(N__16281));
    Odrv4 I__3751 (
            .O(N__16286),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3750 (
            .O(N__16281),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__3749 (
            .O(N__16276),
            .I(N__16273));
    InMux I__3748 (
            .O(N__16273),
            .I(N__16270));
    LocalMux I__3747 (
            .O(N__16270),
            .I(N__16267));
    Span4Mux_h I__3746 (
            .O(N__16267),
            .I(N__16264));
    Odrv4 I__3745 (
            .O(N__16264),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6QZ0));
    InMux I__3744 (
            .O(N__16261),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__3743 (
            .O(N__16258),
            .I(N__16255));
    LocalMux I__3742 (
            .O(N__16255),
            .I(N__16252));
    Span4Mux_h I__3741 (
            .O(N__16252),
            .I(N__16249));
    Odrv4 I__3740 (
            .O(N__16249),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__3739 (
            .O(N__16246),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__3738 (
            .O(N__16243),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__3737 (
            .O(N__16240),
            .I(N__16237));
    LocalMux I__3736 (
            .O(N__16237),
            .I(N__16232));
    InMux I__3735 (
            .O(N__16236),
            .I(N__16229));
    InMux I__3734 (
            .O(N__16235),
            .I(N__16226));
    Span4Mux_v I__3733 (
            .O(N__16232),
            .I(N__16221));
    LocalMux I__3732 (
            .O(N__16229),
            .I(N__16221));
    LocalMux I__3731 (
            .O(N__16226),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0));
    Odrv4 I__3730 (
            .O(N__16221),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0));
    InMux I__3729 (
            .O(N__16216),
            .I(N__16213));
    LocalMux I__3728 (
            .O(N__16213),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0));
    InMux I__3727 (
            .O(N__16210),
            .I(N__16204));
    CascadeMux I__3726 (
            .O(N__16209),
            .I(N__16195));
    CascadeMux I__3725 (
            .O(N__16208),
            .I(N__16192));
    InMux I__3724 (
            .O(N__16207),
            .I(N__16187));
    LocalMux I__3723 (
            .O(N__16204),
            .I(N__16180));
    InMux I__3722 (
            .O(N__16203),
            .I(N__16173));
    InMux I__3721 (
            .O(N__16202),
            .I(N__16173));
    InMux I__3720 (
            .O(N__16201),
            .I(N__16173));
    InMux I__3719 (
            .O(N__16200),
            .I(N__16166));
    InMux I__3718 (
            .O(N__16199),
            .I(N__16166));
    InMux I__3717 (
            .O(N__16198),
            .I(N__16166));
    InMux I__3716 (
            .O(N__16195),
            .I(N__16157));
    InMux I__3715 (
            .O(N__16192),
            .I(N__16157));
    InMux I__3714 (
            .O(N__16191),
            .I(N__16157));
    InMux I__3713 (
            .O(N__16190),
            .I(N__16157));
    LocalMux I__3712 (
            .O(N__16187),
            .I(N__16148));
    InMux I__3711 (
            .O(N__16186),
            .I(N__16139));
    InMux I__3710 (
            .O(N__16185),
            .I(N__16139));
    InMux I__3709 (
            .O(N__16184),
            .I(N__16139));
    InMux I__3708 (
            .O(N__16183),
            .I(N__16139));
    Span4Mux_s2_h I__3707 (
            .O(N__16180),
            .I(N__16129));
    LocalMux I__3706 (
            .O(N__16173),
            .I(N__16129));
    LocalMux I__3705 (
            .O(N__16166),
            .I(N__16129));
    LocalMux I__3704 (
            .O(N__16157),
            .I(N__16129));
    InMux I__3703 (
            .O(N__16156),
            .I(N__16126));
    CascadeMux I__3702 (
            .O(N__16155),
            .I(N__16123));
    InMux I__3701 (
            .O(N__16154),
            .I(N__16120));
    InMux I__3700 (
            .O(N__16153),
            .I(N__16117));
    InMux I__3699 (
            .O(N__16152),
            .I(N__16112));
    InMux I__3698 (
            .O(N__16151),
            .I(N__16112));
    Span4Mux_s3_h I__3697 (
            .O(N__16148),
            .I(N__16107));
    LocalMux I__3696 (
            .O(N__16139),
            .I(N__16107));
    InMux I__3695 (
            .O(N__16138),
            .I(N__16104));
    Span4Mux_h I__3694 (
            .O(N__16129),
            .I(N__16099));
    LocalMux I__3693 (
            .O(N__16126),
            .I(N__16099));
    InMux I__3692 (
            .O(N__16123),
            .I(N__16096));
    LocalMux I__3691 (
            .O(N__16120),
            .I(CO3_0));
    LocalMux I__3690 (
            .O(N__16117),
            .I(CO3_0));
    LocalMux I__3689 (
            .O(N__16112),
            .I(CO3_0));
    Odrv4 I__3688 (
            .O(N__16107),
            .I(CO3_0));
    LocalMux I__3687 (
            .O(N__16104),
            .I(CO3_0));
    Odrv4 I__3686 (
            .O(N__16099),
            .I(CO3_0));
    LocalMux I__3685 (
            .O(N__16096),
            .I(CO3_0));
    InMux I__3684 (
            .O(N__16081),
            .I(N__16078));
    LocalMux I__3683 (
            .O(N__16078),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i));
    InMux I__3682 (
            .O(N__16075),
            .I(N__16063));
    InMux I__3681 (
            .O(N__16074),
            .I(N__16063));
    InMux I__3680 (
            .O(N__16073),
            .I(N__16063));
    InMux I__3679 (
            .O(N__16072),
            .I(N__16063));
    LocalMux I__3678 (
            .O(N__16063),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    CascadeMux I__3677 (
            .O(N__16060),
            .I(N__16057));
    InMux I__3676 (
            .O(N__16057),
            .I(N__16054));
    LocalMux I__3675 (
            .O(N__16054),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKNZ0));
    InMux I__3674 (
            .O(N__16051),
            .I(N__16048));
    LocalMux I__3673 (
            .O(N__16048),
            .I(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5));
    InMux I__3672 (
            .O(N__16045),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__3671 (
            .O(N__16042),
            .I(N__16039));
    LocalMux I__3670 (
            .O(N__16039),
            .I(N__16036));
    Odrv12 I__3669 (
            .O(N__16036),
            .I(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5));
    InMux I__3668 (
            .O(N__16033),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__3667 (
            .O(N__16030),
            .I(N__16025));
    InMux I__3666 (
            .O(N__16029),
            .I(N__15993));
    InMux I__3665 (
            .O(N__16028),
            .I(N__15990));
    InMux I__3664 (
            .O(N__16025),
            .I(N__15985));
    InMux I__3663 (
            .O(N__16024),
            .I(N__15985));
    InMux I__3662 (
            .O(N__16023),
            .I(N__15975));
    InMux I__3661 (
            .O(N__16022),
            .I(N__15975));
    InMux I__3660 (
            .O(N__16021),
            .I(N__15975));
    InMux I__3659 (
            .O(N__16020),
            .I(N__15972));
    InMux I__3658 (
            .O(N__16019),
            .I(N__15965));
    InMux I__3657 (
            .O(N__16018),
            .I(N__15965));
    InMux I__3656 (
            .O(N__16017),
            .I(N__15965));
    InMux I__3655 (
            .O(N__16016),
            .I(N__15962));
    InMux I__3654 (
            .O(N__16015),
            .I(N__15955));
    InMux I__3653 (
            .O(N__16014),
            .I(N__15955));
    InMux I__3652 (
            .O(N__16013),
            .I(N__15955));
    InMux I__3651 (
            .O(N__16012),
            .I(N__15950));
    InMux I__3650 (
            .O(N__16011),
            .I(N__15950));
    InMux I__3649 (
            .O(N__16010),
            .I(N__15945));
    InMux I__3648 (
            .O(N__16009),
            .I(N__15945));
    InMux I__3647 (
            .O(N__16008),
            .I(N__15936));
    InMux I__3646 (
            .O(N__16007),
            .I(N__15936));
    InMux I__3645 (
            .O(N__16006),
            .I(N__15936));
    InMux I__3644 (
            .O(N__16005),
            .I(N__15936));
    InMux I__3643 (
            .O(N__16004),
            .I(N__15927));
    InMux I__3642 (
            .O(N__16003),
            .I(N__15927));
    InMux I__3641 (
            .O(N__16002),
            .I(N__15927));
    InMux I__3640 (
            .O(N__16001),
            .I(N__15927));
    InMux I__3639 (
            .O(N__16000),
            .I(N__15920));
    InMux I__3638 (
            .O(N__15999),
            .I(N__15920));
    InMux I__3637 (
            .O(N__15998),
            .I(N__15920));
    InMux I__3636 (
            .O(N__15997),
            .I(N__15912));
    InMux I__3635 (
            .O(N__15996),
            .I(N__15912));
    LocalMux I__3634 (
            .O(N__15993),
            .I(N__15905));
    LocalMux I__3633 (
            .O(N__15990),
            .I(N__15905));
    LocalMux I__3632 (
            .O(N__15985),
            .I(N__15905));
    InMux I__3631 (
            .O(N__15984),
            .I(N__15898));
    InMux I__3630 (
            .O(N__15983),
            .I(N__15898));
    InMux I__3629 (
            .O(N__15982),
            .I(N__15898));
    LocalMux I__3628 (
            .O(N__15975),
            .I(N__15891));
    LocalMux I__3627 (
            .O(N__15972),
            .I(N__15891));
    LocalMux I__3626 (
            .O(N__15965),
            .I(N__15891));
    LocalMux I__3625 (
            .O(N__15962),
            .I(N__15888));
    LocalMux I__3624 (
            .O(N__15955),
            .I(N__15875));
    LocalMux I__3623 (
            .O(N__15950),
            .I(N__15875));
    LocalMux I__3622 (
            .O(N__15945),
            .I(N__15875));
    LocalMux I__3621 (
            .O(N__15936),
            .I(N__15875));
    LocalMux I__3620 (
            .O(N__15927),
            .I(N__15875));
    LocalMux I__3619 (
            .O(N__15920),
            .I(N__15875));
    InMux I__3618 (
            .O(N__15919),
            .I(N__15870));
    InMux I__3617 (
            .O(N__15918),
            .I(N__15870));
    CascadeMux I__3616 (
            .O(N__15917),
            .I(N__15863));
    LocalMux I__3615 (
            .O(N__15912),
            .I(N__15854));
    Span4Mux_h I__3614 (
            .O(N__15905),
            .I(N__15854));
    LocalMux I__3613 (
            .O(N__15898),
            .I(N__15854));
    Span4Mux_v I__3612 (
            .O(N__15891),
            .I(N__15851));
    Span4Mux_h I__3611 (
            .O(N__15888),
            .I(N__15844));
    Span4Mux_v I__3610 (
            .O(N__15875),
            .I(N__15844));
    LocalMux I__3609 (
            .O(N__15870),
            .I(N__15844));
    InMux I__3608 (
            .O(N__15869),
            .I(N__15841));
    InMux I__3607 (
            .O(N__15868),
            .I(N__15828));
    InMux I__3606 (
            .O(N__15867),
            .I(N__15828));
    InMux I__3605 (
            .O(N__15866),
            .I(N__15828));
    InMux I__3604 (
            .O(N__15863),
            .I(N__15828));
    InMux I__3603 (
            .O(N__15862),
            .I(N__15828));
    InMux I__3602 (
            .O(N__15861),
            .I(N__15828));
    Odrv4 I__3601 (
            .O(N__15854),
            .I(un5_rowlto1));
    Odrv4 I__3600 (
            .O(N__15851),
            .I(un5_rowlto1));
    Odrv4 I__3599 (
            .O(N__15844),
            .I(un5_rowlto1));
    LocalMux I__3598 (
            .O(N__15841),
            .I(un5_rowlto1));
    LocalMux I__3597 (
            .O(N__15828),
            .I(un5_rowlto1));
    CascadeMux I__3596 (
            .O(N__15817),
            .I(N__15809));
    CascadeMux I__3595 (
            .O(N__15816),
            .I(N__15800));
    CascadeMux I__3594 (
            .O(N__15815),
            .I(N__15797));
    InMux I__3593 (
            .O(N__15814),
            .I(N__15784));
    InMux I__3592 (
            .O(N__15813),
            .I(N__15784));
    InMux I__3591 (
            .O(N__15812),
            .I(N__15779));
    InMux I__3590 (
            .O(N__15809),
            .I(N__15779));
    InMux I__3589 (
            .O(N__15808),
            .I(N__15776));
    InMux I__3588 (
            .O(N__15807),
            .I(N__15771));
    InMux I__3587 (
            .O(N__15806),
            .I(N__15771));
    InMux I__3586 (
            .O(N__15805),
            .I(N__15762));
    InMux I__3585 (
            .O(N__15804),
            .I(N__15762));
    InMux I__3584 (
            .O(N__15803),
            .I(N__15762));
    InMux I__3583 (
            .O(N__15800),
            .I(N__15748));
    InMux I__3582 (
            .O(N__15797),
            .I(N__15748));
    InMux I__3581 (
            .O(N__15796),
            .I(N__15737));
    InMux I__3580 (
            .O(N__15795),
            .I(N__15737));
    InMux I__3579 (
            .O(N__15794),
            .I(N__15737));
    InMux I__3578 (
            .O(N__15793),
            .I(N__15737));
    InMux I__3577 (
            .O(N__15792),
            .I(N__15737));
    InMux I__3576 (
            .O(N__15791),
            .I(N__15734));
    InMux I__3575 (
            .O(N__15790),
            .I(N__15729));
    InMux I__3574 (
            .O(N__15789),
            .I(N__15729));
    LocalMux I__3573 (
            .O(N__15784),
            .I(N__15723));
    LocalMux I__3572 (
            .O(N__15779),
            .I(N__15723));
    LocalMux I__3571 (
            .O(N__15776),
            .I(N__15718));
    LocalMux I__3570 (
            .O(N__15771),
            .I(N__15718));
    InMux I__3569 (
            .O(N__15770),
            .I(N__15713));
    InMux I__3568 (
            .O(N__15769),
            .I(N__15713));
    LocalMux I__3567 (
            .O(N__15762),
            .I(N__15710));
    InMux I__3566 (
            .O(N__15761),
            .I(N__15697));
    InMux I__3565 (
            .O(N__15760),
            .I(N__15697));
    InMux I__3564 (
            .O(N__15759),
            .I(N__15697));
    InMux I__3563 (
            .O(N__15758),
            .I(N__15697));
    InMux I__3562 (
            .O(N__15757),
            .I(N__15697));
    InMux I__3561 (
            .O(N__15756),
            .I(N__15697));
    InMux I__3560 (
            .O(N__15755),
            .I(N__15685));
    InMux I__3559 (
            .O(N__15754),
            .I(N__15685));
    InMux I__3558 (
            .O(N__15753),
            .I(N__15685));
    LocalMux I__3557 (
            .O(N__15748),
            .I(N__15677));
    LocalMux I__3556 (
            .O(N__15737),
            .I(N__15677));
    LocalMux I__3555 (
            .O(N__15734),
            .I(N__15677));
    LocalMux I__3554 (
            .O(N__15729),
            .I(N__15674));
    InMux I__3553 (
            .O(N__15728),
            .I(N__15671));
    Span4Mux_v I__3552 (
            .O(N__15723),
            .I(N__15664));
    Span4Mux_v I__3551 (
            .O(N__15718),
            .I(N__15664));
    LocalMux I__3550 (
            .O(N__15713),
            .I(N__15664));
    Span4Mux_v I__3549 (
            .O(N__15710),
            .I(N__15659));
    LocalMux I__3548 (
            .O(N__15697),
            .I(N__15659));
    InMux I__3547 (
            .O(N__15696),
            .I(N__15648));
    InMux I__3546 (
            .O(N__15695),
            .I(N__15648));
    InMux I__3545 (
            .O(N__15694),
            .I(N__15648));
    InMux I__3544 (
            .O(N__15693),
            .I(N__15648));
    InMux I__3543 (
            .O(N__15692),
            .I(N__15648));
    LocalMux I__3542 (
            .O(N__15685),
            .I(N__15645));
    InMux I__3541 (
            .O(N__15684),
            .I(N__15642));
    Span4Mux_h I__3540 (
            .O(N__15677),
            .I(N__15639));
    Odrv4 I__3539 (
            .O(N__15674),
            .I(un5_rowlto0));
    LocalMux I__3538 (
            .O(N__15671),
            .I(un5_rowlto0));
    Odrv4 I__3537 (
            .O(N__15664),
            .I(un5_rowlto0));
    Odrv4 I__3536 (
            .O(N__15659),
            .I(un5_rowlto0));
    LocalMux I__3535 (
            .O(N__15648),
            .I(un5_rowlto0));
    Odrv12 I__3534 (
            .O(N__15645),
            .I(un5_rowlto0));
    LocalMux I__3533 (
            .O(N__15642),
            .I(un5_rowlto0));
    Odrv4 I__3532 (
            .O(N__15639),
            .I(un5_rowlto0));
    CascadeMux I__3531 (
            .O(N__15622),
            .I(un5_rowlto1_cascade_));
    CascadeMux I__3530 (
            .O(N__15619),
            .I(N__15613));
    CascadeMux I__3529 (
            .O(N__15618),
            .I(N__15610));
    InMux I__3528 (
            .O(N__15617),
            .I(N__15605));
    InMux I__3527 (
            .O(N__15616),
            .I(N__15602));
    InMux I__3526 (
            .O(N__15613),
            .I(N__15595));
    InMux I__3525 (
            .O(N__15610),
            .I(N__15595));
    InMux I__3524 (
            .O(N__15609),
            .I(N__15595));
    InMux I__3523 (
            .O(N__15608),
            .I(N__15581));
    LocalMux I__3522 (
            .O(N__15605),
            .I(N__15574));
    LocalMux I__3521 (
            .O(N__15602),
            .I(N__15571));
    LocalMux I__3520 (
            .O(N__15595),
            .I(N__15568));
    InMux I__3519 (
            .O(N__15594),
            .I(N__15563));
    InMux I__3518 (
            .O(N__15593),
            .I(N__15563));
    InMux I__3517 (
            .O(N__15592),
            .I(N__15560));
    InMux I__3516 (
            .O(N__15591),
            .I(N__15555));
    InMux I__3515 (
            .O(N__15590),
            .I(N__15555));
    InMux I__3514 (
            .O(N__15589),
            .I(N__15552));
    InMux I__3513 (
            .O(N__15588),
            .I(N__15549));
    InMux I__3512 (
            .O(N__15587),
            .I(N__15546));
    InMux I__3511 (
            .O(N__15586),
            .I(N__15541));
    InMux I__3510 (
            .O(N__15585),
            .I(N__15538));
    InMux I__3509 (
            .O(N__15584),
            .I(N__15535));
    LocalMux I__3508 (
            .O(N__15581),
            .I(N__15532));
    InMux I__3507 (
            .O(N__15580),
            .I(N__15529));
    InMux I__3506 (
            .O(N__15579),
            .I(N__15526));
    InMux I__3505 (
            .O(N__15578),
            .I(N__15521));
    InMux I__3504 (
            .O(N__15577),
            .I(N__15521));
    Span4Mux_s1_h I__3503 (
            .O(N__15574),
            .I(N__15512));
    Span4Mux_v I__3502 (
            .O(N__15571),
            .I(N__15512));
    Span4Mux_v I__3501 (
            .O(N__15568),
            .I(N__15512));
    LocalMux I__3500 (
            .O(N__15563),
            .I(N__15512));
    LocalMux I__3499 (
            .O(N__15560),
            .I(N__15505));
    LocalMux I__3498 (
            .O(N__15555),
            .I(N__15505));
    LocalMux I__3497 (
            .O(N__15552),
            .I(N__15505));
    LocalMux I__3496 (
            .O(N__15549),
            .I(N__15500));
    LocalMux I__3495 (
            .O(N__15546),
            .I(N__15500));
    CascadeMux I__3494 (
            .O(N__15545),
            .I(N__15496));
    CascadeMux I__3493 (
            .O(N__15544),
            .I(N__15493));
    LocalMux I__3492 (
            .O(N__15541),
            .I(N__15489));
    LocalMux I__3491 (
            .O(N__15538),
            .I(N__15486));
    LocalMux I__3490 (
            .O(N__15535),
            .I(N__15475));
    Span4Mux_h I__3489 (
            .O(N__15532),
            .I(N__15475));
    LocalMux I__3488 (
            .O(N__15529),
            .I(N__15475));
    LocalMux I__3487 (
            .O(N__15526),
            .I(N__15475));
    LocalMux I__3486 (
            .O(N__15521),
            .I(N__15475));
    Span4Mux_h I__3485 (
            .O(N__15512),
            .I(N__15472));
    Span4Mux_v I__3484 (
            .O(N__15505),
            .I(N__15467));
    Span4Mux_h I__3483 (
            .O(N__15500),
            .I(N__15467));
    InMux I__3482 (
            .O(N__15499),
            .I(N__15464));
    InMux I__3481 (
            .O(N__15496),
            .I(N__15457));
    InMux I__3480 (
            .O(N__15493),
            .I(N__15457));
    InMux I__3479 (
            .O(N__15492),
            .I(N__15457));
    Odrv4 I__3478 (
            .O(N__15489),
            .I(un5_rowlto3));
    Odrv12 I__3477 (
            .O(N__15486),
            .I(un5_rowlto3));
    Odrv4 I__3476 (
            .O(N__15475),
            .I(un5_rowlto3));
    Odrv4 I__3475 (
            .O(N__15472),
            .I(un5_rowlto3));
    Odrv4 I__3474 (
            .O(N__15467),
            .I(un5_rowlto3));
    LocalMux I__3473 (
            .O(N__15464),
            .I(un5_rowlto3));
    LocalMux I__3472 (
            .O(N__15457),
            .I(un5_rowlto3));
    InMux I__3471 (
            .O(N__15442),
            .I(N__15439));
    LocalMux I__3470 (
            .O(N__15439),
            .I(N__15436));
    Span4Mux_h I__3469 (
            .O(N__15436),
            .I(N__15433));
    Odrv4 I__3468 (
            .O(N__15433),
            .I(un116_pixel_2_am_0));
    CascadeMux I__3467 (
            .O(N__15430),
            .I(N__15426));
    InMux I__3466 (
            .O(N__15429),
            .I(N__15421));
    InMux I__3465 (
            .O(N__15426),
            .I(N__15421));
    LocalMux I__3464 (
            .O(N__15421),
            .I(N__15418));
    Span4Mux_s1_h I__3463 (
            .O(N__15418),
            .I(N__15415));
    Odrv4 I__3462 (
            .O(N__15415),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    InMux I__3461 (
            .O(N__15412),
            .I(N__15409));
    LocalMux I__3460 (
            .O(N__15409),
            .I(if_generate_plus_mult1_un75_sum_axb_4_l_fx));
    CascadeMux I__3459 (
            .O(N__15406),
            .I(N__15390));
    CascadeMux I__3458 (
            .O(N__15405),
            .I(N__15386));
    CascadeMux I__3457 (
            .O(N__15404),
            .I(N__15377));
    InMux I__3456 (
            .O(N__15403),
            .I(N__15368));
    InMux I__3455 (
            .O(N__15402),
            .I(N__15368));
    InMux I__3454 (
            .O(N__15401),
            .I(N__15368));
    InMux I__3453 (
            .O(N__15400),
            .I(N__15357));
    InMux I__3452 (
            .O(N__15399),
            .I(N__15357));
    InMux I__3451 (
            .O(N__15398),
            .I(N__15357));
    InMux I__3450 (
            .O(N__15397),
            .I(N__15357));
    InMux I__3449 (
            .O(N__15396),
            .I(N__15357));
    InMux I__3448 (
            .O(N__15395),
            .I(N__15349));
    InMux I__3447 (
            .O(N__15394),
            .I(N__15349));
    InMux I__3446 (
            .O(N__15393),
            .I(N__15338));
    InMux I__3445 (
            .O(N__15390),
            .I(N__15338));
    InMux I__3444 (
            .O(N__15389),
            .I(N__15338));
    InMux I__3443 (
            .O(N__15386),
            .I(N__15338));
    InMux I__3442 (
            .O(N__15385),
            .I(N__15338));
    CascadeMux I__3441 (
            .O(N__15384),
            .I(N__15330));
    CascadeMux I__3440 (
            .O(N__15383),
            .I(N__15327));
    InMux I__3439 (
            .O(N__15382),
            .I(N__15323));
    InMux I__3438 (
            .O(N__15381),
            .I(N__15312));
    InMux I__3437 (
            .O(N__15380),
            .I(N__15312));
    InMux I__3436 (
            .O(N__15377),
            .I(N__15312));
    InMux I__3435 (
            .O(N__15376),
            .I(N__15312));
    InMux I__3434 (
            .O(N__15375),
            .I(N__15312));
    LocalMux I__3433 (
            .O(N__15368),
            .I(N__15309));
    LocalMux I__3432 (
            .O(N__15357),
            .I(N__15306));
    InMux I__3431 (
            .O(N__15356),
            .I(N__15303));
    InMux I__3430 (
            .O(N__15355),
            .I(N__15289));
    InMux I__3429 (
            .O(N__15354),
            .I(N__15289));
    LocalMux I__3428 (
            .O(N__15349),
            .I(N__15282));
    LocalMux I__3427 (
            .O(N__15338),
            .I(N__15282));
    InMux I__3426 (
            .O(N__15337),
            .I(N__15277));
    InMux I__3425 (
            .O(N__15336),
            .I(N__15277));
    InMux I__3424 (
            .O(N__15335),
            .I(N__15272));
    InMux I__3423 (
            .O(N__15334),
            .I(N__15272));
    InMux I__3422 (
            .O(N__15333),
            .I(N__15269));
    InMux I__3421 (
            .O(N__15330),
            .I(N__15262));
    InMux I__3420 (
            .O(N__15327),
            .I(N__15262));
    InMux I__3419 (
            .O(N__15326),
            .I(N__15262));
    LocalMux I__3418 (
            .O(N__15323),
            .I(N__15259));
    LocalMux I__3417 (
            .O(N__15312),
            .I(N__15250));
    Span4Mux_v I__3416 (
            .O(N__15309),
            .I(N__15250));
    Span4Mux_v I__3415 (
            .O(N__15306),
            .I(N__15250));
    LocalMux I__3414 (
            .O(N__15303),
            .I(N__15250));
    InMux I__3413 (
            .O(N__15302),
            .I(N__15244));
    InMux I__3412 (
            .O(N__15301),
            .I(N__15244));
    InMux I__3411 (
            .O(N__15300),
            .I(N__15241));
    InMux I__3410 (
            .O(N__15299),
            .I(N__15234));
    InMux I__3409 (
            .O(N__15298),
            .I(N__15234));
    InMux I__3408 (
            .O(N__15297),
            .I(N__15234));
    InMux I__3407 (
            .O(N__15296),
            .I(N__15229));
    InMux I__3406 (
            .O(N__15295),
            .I(N__15229));
    InMux I__3405 (
            .O(N__15294),
            .I(N__15226));
    LocalMux I__3404 (
            .O(N__15289),
            .I(N__15223));
    InMux I__3403 (
            .O(N__15288),
            .I(N__15220));
    InMux I__3402 (
            .O(N__15287),
            .I(N__15217));
    Span4Mux_v I__3401 (
            .O(N__15282),
            .I(N__15214));
    LocalMux I__3400 (
            .O(N__15277),
            .I(N__15205));
    LocalMux I__3399 (
            .O(N__15272),
            .I(N__15205));
    LocalMux I__3398 (
            .O(N__15269),
            .I(N__15205));
    LocalMux I__3397 (
            .O(N__15262),
            .I(N__15205));
    Span4Mux_v I__3396 (
            .O(N__15259),
            .I(N__15200));
    Span4Mux_h I__3395 (
            .O(N__15250),
            .I(N__15200));
    InMux I__3394 (
            .O(N__15249),
            .I(N__15197));
    LocalMux I__3393 (
            .O(N__15244),
            .I(N__15190));
    LocalMux I__3392 (
            .O(N__15241),
            .I(N__15190));
    LocalMux I__3391 (
            .O(N__15234),
            .I(N__15190));
    LocalMux I__3390 (
            .O(N__15229),
            .I(un5_rowlto2));
    LocalMux I__3389 (
            .O(N__15226),
            .I(un5_rowlto2));
    Odrv12 I__3388 (
            .O(N__15223),
            .I(un5_rowlto2));
    LocalMux I__3387 (
            .O(N__15220),
            .I(un5_rowlto2));
    LocalMux I__3386 (
            .O(N__15217),
            .I(un5_rowlto2));
    Odrv4 I__3385 (
            .O(N__15214),
            .I(un5_rowlto2));
    Odrv4 I__3384 (
            .O(N__15205),
            .I(un5_rowlto2));
    Odrv4 I__3383 (
            .O(N__15200),
            .I(un5_rowlto2));
    LocalMux I__3382 (
            .O(N__15197),
            .I(un5_rowlto2));
    Odrv12 I__3381 (
            .O(N__15190),
            .I(un5_rowlto2));
    InMux I__3380 (
            .O(N__15169),
            .I(N__15166));
    LocalMux I__3379 (
            .O(N__15166),
            .I(un5_rowlto2_i));
    InMux I__3378 (
            .O(N__15163),
            .I(N__15159));
    InMux I__3377 (
            .O(N__15162),
            .I(N__15156));
    LocalMux I__3376 (
            .O(N__15159),
            .I(N__15152));
    LocalMux I__3375 (
            .O(N__15156),
            .I(N__15149));
    InMux I__3374 (
            .O(N__15155),
            .I(N__15145));
    Span4Mux_v I__3373 (
            .O(N__15152),
            .I(N__15140));
    Span4Mux_s1_h I__3372 (
            .O(N__15149),
            .I(N__15140));
    InMux I__3371 (
            .O(N__15148),
            .I(N__15137));
    LocalMux I__3370 (
            .O(N__15145),
            .I(N__15134));
    Span4Mux_h I__3369 (
            .O(N__15140),
            .I(N__15131));
    LocalMux I__3368 (
            .O(N__15137),
            .I(N__15126));
    Span4Mux_v I__3367 (
            .O(N__15134),
            .I(N__15126));
    Odrv4 I__3366 (
            .O(N__15131),
            .I(charx_if_generate_plus_mult1_un68_sum));
    Odrv4 I__3365 (
            .O(N__15126),
            .I(charx_if_generate_plus_mult1_un68_sum));
    CascadeMux I__3364 (
            .O(N__15121),
            .I(N__15118));
    InMux I__3363 (
            .O(N__15118),
            .I(N__15115));
    LocalMux I__3362 (
            .O(N__15115),
            .I(N__15112));
    Odrv4 I__3361 (
            .O(N__15112),
            .I(column_1_if_generate_plus_mult1_un75_sum_iZ0));
    InMux I__3360 (
            .O(N__15109),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    CascadeMux I__3359 (
            .O(N__15106),
            .I(N__15103));
    InMux I__3358 (
            .O(N__15103),
            .I(N__15099));
    InMux I__3357 (
            .O(N__15102),
            .I(N__15094));
    LocalMux I__3356 (
            .O(N__15099),
            .I(N__15090));
    InMux I__3355 (
            .O(N__15098),
            .I(N__15085));
    InMux I__3354 (
            .O(N__15097),
            .I(N__15085));
    LocalMux I__3353 (
            .O(N__15094),
            .I(N__15082));
    CascadeMux I__3352 (
            .O(N__15093),
            .I(N__15078));
    Span4Mux_v I__3351 (
            .O(N__15090),
            .I(N__15072));
    LocalMux I__3350 (
            .O(N__15085),
            .I(N__15072));
    Span4Mux_s1_h I__3349 (
            .O(N__15082),
            .I(N__15069));
    InMux I__3348 (
            .O(N__15081),
            .I(N__15066));
    InMux I__3347 (
            .O(N__15078),
            .I(N__15062));
    InMux I__3346 (
            .O(N__15077),
            .I(N__15059));
    Span4Mux_h I__3345 (
            .O(N__15072),
            .I(N__15056));
    Span4Mux_h I__3344 (
            .O(N__15069),
            .I(N__15051));
    LocalMux I__3343 (
            .O(N__15066),
            .I(N__15051));
    InMux I__3342 (
            .O(N__15065),
            .I(N__15048));
    LocalMux I__3341 (
            .O(N__15062),
            .I(N__15045));
    LocalMux I__3340 (
            .O(N__15059),
            .I(charx_if_generate_plus_mult1_un26_sum));
    Odrv4 I__3339 (
            .O(N__15056),
            .I(charx_if_generate_plus_mult1_un26_sum));
    Odrv4 I__3338 (
            .O(N__15051),
            .I(charx_if_generate_plus_mult1_un26_sum));
    LocalMux I__3337 (
            .O(N__15048),
            .I(charx_if_generate_plus_mult1_un26_sum));
    Odrv4 I__3336 (
            .O(N__15045),
            .I(charx_if_generate_plus_mult1_un26_sum));
    InMux I__3335 (
            .O(N__15034),
            .I(N__15031));
    LocalMux I__3334 (
            .O(N__15031),
            .I(G_346));
    InMux I__3333 (
            .O(N__15028),
            .I(column_1_if_generate_plus_mult1_un82_sum_cry_4));
    CascadeMux I__3332 (
            .O(N__15025),
            .I(un5_rowlto0_cascade_));
    InMux I__3331 (
            .O(N__15022),
            .I(N__15019));
    LocalMux I__3330 (
            .O(N__15019),
            .I(un116_pixel_1_bmZ0Z_1));
    CascadeMux I__3329 (
            .O(N__15016),
            .I(N__15004));
    CascadeMux I__3328 (
            .O(N__15015),
            .I(N__15000));
    CascadeMux I__3327 (
            .O(N__15014),
            .I(N__14996));
    InMux I__3326 (
            .O(N__15013),
            .I(N__14991));
    CascadeMux I__3325 (
            .O(N__15012),
            .I(N__14988));
    InMux I__3324 (
            .O(N__15011),
            .I(N__14977));
    InMux I__3323 (
            .O(N__15010),
            .I(N__14977));
    InMux I__3322 (
            .O(N__15009),
            .I(N__14977));
    CascadeMux I__3321 (
            .O(N__15008),
            .I(N__14971));
    InMux I__3320 (
            .O(N__15007),
            .I(N__14968));
    InMux I__3319 (
            .O(N__15004),
            .I(N__14965));
    InMux I__3318 (
            .O(N__15003),
            .I(N__14960));
    InMux I__3317 (
            .O(N__15000),
            .I(N__14960));
    InMux I__3316 (
            .O(N__14999),
            .I(N__14955));
    InMux I__3315 (
            .O(N__14996),
            .I(N__14955));
    CascadeMux I__3314 (
            .O(N__14995),
            .I(N__14951));
    InMux I__3313 (
            .O(N__14994),
            .I(N__14946));
    LocalMux I__3312 (
            .O(N__14991),
            .I(N__14943));
    InMux I__3311 (
            .O(N__14988),
            .I(N__14940));
    InMux I__3310 (
            .O(N__14987),
            .I(N__14935));
    InMux I__3309 (
            .O(N__14986),
            .I(N__14935));
    InMux I__3308 (
            .O(N__14985),
            .I(N__14930));
    InMux I__3307 (
            .O(N__14984),
            .I(N__14930));
    LocalMux I__3306 (
            .O(N__14977),
            .I(N__14927));
    CascadeMux I__3305 (
            .O(N__14976),
            .I(N__14924));
    CascadeMux I__3304 (
            .O(N__14975),
            .I(N__14921));
    InMux I__3303 (
            .O(N__14974),
            .I(N__14917));
    InMux I__3302 (
            .O(N__14971),
            .I(N__14914));
    LocalMux I__3301 (
            .O(N__14968),
            .I(N__14909));
    LocalMux I__3300 (
            .O(N__14965),
            .I(N__14909));
    LocalMux I__3299 (
            .O(N__14960),
            .I(N__14904));
    LocalMux I__3298 (
            .O(N__14955),
            .I(N__14904));
    InMux I__3297 (
            .O(N__14954),
            .I(N__14897));
    InMux I__3296 (
            .O(N__14951),
            .I(N__14894));
    InMux I__3295 (
            .O(N__14950),
            .I(N__14889));
    InMux I__3294 (
            .O(N__14949),
            .I(N__14889));
    LocalMux I__3293 (
            .O(N__14946),
            .I(N__14886));
    Span4Mux_s2_h I__3292 (
            .O(N__14943),
            .I(N__14883));
    LocalMux I__3291 (
            .O(N__14940),
            .I(N__14874));
    LocalMux I__3290 (
            .O(N__14935),
            .I(N__14874));
    LocalMux I__3289 (
            .O(N__14930),
            .I(N__14874));
    Span4Mux_s1_h I__3288 (
            .O(N__14927),
            .I(N__14874));
    InMux I__3287 (
            .O(N__14924),
            .I(N__14871));
    InMux I__3286 (
            .O(N__14921),
            .I(N__14868));
    InMux I__3285 (
            .O(N__14920),
            .I(N__14865));
    LocalMux I__3284 (
            .O(N__14917),
            .I(N__14862));
    LocalMux I__3283 (
            .O(N__14914),
            .I(N__14859));
    Span4Mux_h I__3282 (
            .O(N__14909),
            .I(N__14856));
    Span4Mux_h I__3281 (
            .O(N__14904),
            .I(N__14853));
    InMux I__3280 (
            .O(N__14903),
            .I(N__14850));
    InMux I__3279 (
            .O(N__14902),
            .I(N__14843));
    InMux I__3278 (
            .O(N__14901),
            .I(N__14843));
    InMux I__3277 (
            .O(N__14900),
            .I(N__14843));
    LocalMux I__3276 (
            .O(N__14897),
            .I(N__14836));
    LocalMux I__3275 (
            .O(N__14894),
            .I(N__14836));
    LocalMux I__3274 (
            .O(N__14889),
            .I(N__14836));
    Span4Mux_h I__3273 (
            .O(N__14886),
            .I(N__14829));
    Span4Mux_h I__3272 (
            .O(N__14883),
            .I(N__14829));
    Span4Mux_h I__3271 (
            .O(N__14874),
            .I(N__14829));
    LocalMux I__3270 (
            .O(N__14871),
            .I(N__14822));
    LocalMux I__3269 (
            .O(N__14868),
            .I(N__14822));
    LocalMux I__3268 (
            .O(N__14865),
            .I(N__14822));
    Odrv4 I__3267 (
            .O(N__14862),
            .I(beamYZ0Z_1));
    Odrv12 I__3266 (
            .O(N__14859),
            .I(beamYZ0Z_1));
    Odrv4 I__3265 (
            .O(N__14856),
            .I(beamYZ0Z_1));
    Odrv4 I__3264 (
            .O(N__14853),
            .I(beamYZ0Z_1));
    LocalMux I__3263 (
            .O(N__14850),
            .I(beamYZ0Z_1));
    LocalMux I__3262 (
            .O(N__14843),
            .I(beamYZ0Z_1));
    Odrv12 I__3261 (
            .O(N__14836),
            .I(beamYZ0Z_1));
    Odrv4 I__3260 (
            .O(N__14829),
            .I(beamYZ0Z_1));
    Odrv12 I__3259 (
            .O(N__14822),
            .I(beamYZ0Z_1));
    CascadeMux I__3258 (
            .O(N__14803),
            .I(un116_pixel_1_bmZ0Z_1_cascade_));
    InMux I__3257 (
            .O(N__14800),
            .I(N__14797));
    LocalMux I__3256 (
            .O(N__14797),
            .I(N__14794));
    Span4Mux_h I__3255 (
            .O(N__14794),
            .I(N__14791));
    Odrv4 I__3254 (
            .O(N__14791),
            .I(beamY_RNIV622TRZ0Z_1));
    InMux I__3253 (
            .O(N__14788),
            .I(N__14785));
    LocalMux I__3252 (
            .O(N__14785),
            .I(N__14782));
    Odrv4 I__3251 (
            .O(N__14782),
            .I(un116_pixel_2_ns_1_4));
    CascadeMux I__3250 (
            .O(N__14779),
            .I(N__14770));
    CascadeMux I__3249 (
            .O(N__14778),
            .I(N__14762));
    CascadeMux I__3248 (
            .O(N__14777),
            .I(N__14754));
    CascadeMux I__3247 (
            .O(N__14776),
            .I(N__14747));
    CascadeMux I__3246 (
            .O(N__14775),
            .I(N__14738));
    CascadeMux I__3245 (
            .O(N__14774),
            .I(N__14733));
    CascadeMux I__3244 (
            .O(N__14773),
            .I(N__14730));
    InMux I__3243 (
            .O(N__14770),
            .I(N__14726));
    InMux I__3242 (
            .O(N__14769),
            .I(N__14723));
    InMux I__3241 (
            .O(N__14768),
            .I(N__14714));
    InMux I__3240 (
            .O(N__14767),
            .I(N__14714));
    InMux I__3239 (
            .O(N__14766),
            .I(N__14714));
    InMux I__3238 (
            .O(N__14765),
            .I(N__14714));
    InMux I__3237 (
            .O(N__14762),
            .I(N__14709));
    InMux I__3236 (
            .O(N__14761),
            .I(N__14709));
    InMux I__3235 (
            .O(N__14760),
            .I(N__14706));
    CascadeMux I__3234 (
            .O(N__14759),
            .I(N__14703));
    InMux I__3233 (
            .O(N__14758),
            .I(N__14695));
    InMux I__3232 (
            .O(N__14757),
            .I(N__14695));
    InMux I__3231 (
            .O(N__14754),
            .I(N__14695));
    InMux I__3230 (
            .O(N__14753),
            .I(N__14690));
    InMux I__3229 (
            .O(N__14752),
            .I(N__14690));
    InMux I__3228 (
            .O(N__14751),
            .I(N__14687));
    InMux I__3227 (
            .O(N__14750),
            .I(N__14684));
    InMux I__3226 (
            .O(N__14747),
            .I(N__14681));
    InMux I__3225 (
            .O(N__14746),
            .I(N__14676));
    InMux I__3224 (
            .O(N__14745),
            .I(N__14676));
    CascadeMux I__3223 (
            .O(N__14744),
            .I(N__14673));
    InMux I__3222 (
            .O(N__14743),
            .I(N__14666));
    InMux I__3221 (
            .O(N__14742),
            .I(N__14666));
    InMux I__3220 (
            .O(N__14741),
            .I(N__14666));
    InMux I__3219 (
            .O(N__14738),
            .I(N__14657));
    InMux I__3218 (
            .O(N__14737),
            .I(N__14657));
    InMux I__3217 (
            .O(N__14736),
            .I(N__14657));
    InMux I__3216 (
            .O(N__14733),
            .I(N__14657));
    InMux I__3215 (
            .O(N__14730),
            .I(N__14652));
    InMux I__3214 (
            .O(N__14729),
            .I(N__14652));
    LocalMux I__3213 (
            .O(N__14726),
            .I(N__14645));
    LocalMux I__3212 (
            .O(N__14723),
            .I(N__14645));
    LocalMux I__3211 (
            .O(N__14714),
            .I(N__14645));
    LocalMux I__3210 (
            .O(N__14709),
            .I(N__14642));
    LocalMux I__3209 (
            .O(N__14706),
            .I(N__14638));
    InMux I__3208 (
            .O(N__14703),
            .I(N__14635));
    CascadeMux I__3207 (
            .O(N__14702),
            .I(N__14631));
    LocalMux I__3206 (
            .O(N__14695),
            .I(N__14627));
    LocalMux I__3205 (
            .O(N__14690),
            .I(N__14622));
    LocalMux I__3204 (
            .O(N__14687),
            .I(N__14622));
    LocalMux I__3203 (
            .O(N__14684),
            .I(N__14617));
    LocalMux I__3202 (
            .O(N__14681),
            .I(N__14617));
    LocalMux I__3201 (
            .O(N__14676),
            .I(N__14614));
    InMux I__3200 (
            .O(N__14673),
            .I(N__14611));
    LocalMux I__3199 (
            .O(N__14666),
            .I(N__14608));
    LocalMux I__3198 (
            .O(N__14657),
            .I(N__14599));
    LocalMux I__3197 (
            .O(N__14652),
            .I(N__14599));
    Span4Mux_v I__3196 (
            .O(N__14645),
            .I(N__14599));
    Span4Mux_s1_h I__3195 (
            .O(N__14642),
            .I(N__14599));
    InMux I__3194 (
            .O(N__14641),
            .I(N__14596));
    Span12Mux_s5_h I__3193 (
            .O(N__14638),
            .I(N__14593));
    LocalMux I__3192 (
            .O(N__14635),
            .I(N__14590));
    InMux I__3191 (
            .O(N__14634),
            .I(N__14587));
    InMux I__3190 (
            .O(N__14631),
            .I(N__14582));
    InMux I__3189 (
            .O(N__14630),
            .I(N__14582));
    Span4Mux_h I__3188 (
            .O(N__14627),
            .I(N__14577));
    Span4Mux_h I__3187 (
            .O(N__14622),
            .I(N__14577));
    Span4Mux_h I__3186 (
            .O(N__14617),
            .I(N__14574));
    Span4Mux_v I__3185 (
            .O(N__14614),
            .I(N__14569));
    LocalMux I__3184 (
            .O(N__14611),
            .I(N__14569));
    Span4Mux_v I__3183 (
            .O(N__14608),
            .I(N__14564));
    Span4Mux_h I__3182 (
            .O(N__14599),
            .I(N__14564));
    LocalMux I__3181 (
            .O(N__14596),
            .I(beamYZ0Z_0));
    Odrv12 I__3180 (
            .O(N__14593),
            .I(beamYZ0Z_0));
    Odrv4 I__3179 (
            .O(N__14590),
            .I(beamYZ0Z_0));
    LocalMux I__3178 (
            .O(N__14587),
            .I(beamYZ0Z_0));
    LocalMux I__3177 (
            .O(N__14582),
            .I(beamYZ0Z_0));
    Odrv4 I__3176 (
            .O(N__14577),
            .I(beamYZ0Z_0));
    Odrv4 I__3175 (
            .O(N__14574),
            .I(beamYZ0Z_0));
    Odrv4 I__3174 (
            .O(N__14569),
            .I(beamYZ0Z_0));
    Odrv4 I__3173 (
            .O(N__14564),
            .I(beamYZ0Z_0));
    InMux I__3172 (
            .O(N__14545),
            .I(N__14542));
    LocalMux I__3171 (
            .O(N__14542),
            .I(N__14539));
    Odrv4 I__3170 (
            .O(N__14539),
            .I(beamY_RNIITCG3J3Z0Z_0));
    CascadeMux I__3169 (
            .O(N__14536),
            .I(N__14533));
    InMux I__3168 (
            .O(N__14533),
            .I(N__14530));
    LocalMux I__3167 (
            .O(N__14530),
            .I(N__14527));
    Odrv4 I__3166 (
            .O(N__14527),
            .I(column_1_if_generate_plus_mult1_un68_sum_iZ0));
    InMux I__3165 (
            .O(N__14524),
            .I(N__14521));
    LocalMux I__3164 (
            .O(N__14521),
            .I(if_generate_plus_mult1_un75_sum_cry_2_s));
    InMux I__3163 (
            .O(N__14518),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_1));
    CascadeMux I__3162 (
            .O(N__14515),
            .I(N__14512));
    InMux I__3161 (
            .O(N__14512),
            .I(N__14509));
    LocalMux I__3160 (
            .O(N__14509),
            .I(N__14506));
    Odrv12 I__3159 (
            .O(N__14506),
            .I(if_generate_plus_mult1_un68_sum_cry_2_s));
    CascadeMux I__3158 (
            .O(N__14503),
            .I(N__14500));
    InMux I__3157 (
            .O(N__14500),
            .I(N__14497));
    LocalMux I__3156 (
            .O(N__14497),
            .I(if_generate_plus_mult1_un75_sum_cry_3_s));
    InMux I__3155 (
            .O(N__14494),
            .I(column_1_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__3154 (
            .O(N__14491),
            .I(N__14488));
    LocalMux I__3153 (
            .O(N__14488),
            .I(un116_pixel_2_bmZ0Z_5));
    CascadeMux I__3152 (
            .O(N__14485),
            .I(un114_pixel_7_1_7__N_9_cascade_));
    CascadeMux I__3151 (
            .O(N__14482),
            .I(un114_pixel_1_0_3__un116_pixel_3_ns_1Z0Z_0_cascade_));
    InMux I__3150 (
            .O(N__14479),
            .I(N__14476));
    LocalMux I__3149 (
            .O(N__14476),
            .I(un114_pixel_6_1_5__N_8));
    InMux I__3148 (
            .O(N__14473),
            .I(N__14470));
    LocalMux I__3147 (
            .O(N__14470),
            .I(N__14467));
    Span4Mux_h I__3146 (
            .O(N__14467),
            .I(N__14464));
    Odrv4 I__3145 (
            .O(N__14464),
            .I(N_371));
    InMux I__3144 (
            .O(N__14461),
            .I(N__14458));
    LocalMux I__3143 (
            .O(N__14458),
            .I(N__14455));
    Odrv4 I__3142 (
            .O(N__14455),
            .I(beamY_RNIJUCG3J3Z0Z_1));
    InMux I__3141 (
            .O(N__14452),
            .I(N__14447));
    InMux I__3140 (
            .O(N__14451),
            .I(N__14441));
    InMux I__3139 (
            .O(N__14450),
            .I(N__14438));
    LocalMux I__3138 (
            .O(N__14447),
            .I(N__14435));
    InMux I__3137 (
            .O(N__14446),
            .I(N__14430));
    InMux I__3136 (
            .O(N__14445),
            .I(N__14430));
    InMux I__3135 (
            .O(N__14444),
            .I(N__14427));
    LocalMux I__3134 (
            .O(N__14441),
            .I(N__14420));
    LocalMux I__3133 (
            .O(N__14438),
            .I(N__14420));
    Span4Mux_s3_h I__3132 (
            .O(N__14435),
            .I(N__14415));
    LocalMux I__3131 (
            .O(N__14430),
            .I(N__14415));
    LocalMux I__3130 (
            .O(N__14427),
            .I(N__14412));
    InMux I__3129 (
            .O(N__14426),
            .I(N__14407));
    InMux I__3128 (
            .O(N__14425),
            .I(N__14407));
    Span4Mux_v I__3127 (
            .O(N__14420),
            .I(N__14398));
    Span4Mux_v I__3126 (
            .O(N__14415),
            .I(N__14398));
    Span4Mux_s3_h I__3125 (
            .O(N__14412),
            .I(N__14398));
    LocalMux I__3124 (
            .O(N__14407),
            .I(N__14398));
    Odrv4 I__3123 (
            .O(N__14398),
            .I(charx_if_generate_plus_mult1_un75_sum));
    InMux I__3122 (
            .O(N__14395),
            .I(N__14392));
    LocalMux I__3121 (
            .O(N__14392),
            .I(G_345));
    InMux I__3120 (
            .O(N__14389),
            .I(N__14383));
    InMux I__3119 (
            .O(N__14388),
            .I(N__14383));
    LocalMux I__3118 (
            .O(N__14383),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8));
    InMux I__3117 (
            .O(N__14380),
            .I(N__14377));
    LocalMux I__3116 (
            .O(N__14377),
            .I(N__14374));
    Odrv4 I__3115 (
            .O(N__14374),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__3114 (
            .O(N__14371),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__3113 (
            .O(N__14368),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7));
    InMux I__3112 (
            .O(N__14365),
            .I(N__14362));
    LocalMux I__3111 (
            .O(N__14362),
            .I(N__14357));
    InMux I__3110 (
            .O(N__14361),
            .I(N__14354));
    InMux I__3109 (
            .O(N__14360),
            .I(N__14351));
    Odrv4 I__3108 (
            .O(N__14357),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052));
    LocalMux I__3107 (
            .O(N__14354),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052));
    LocalMux I__3106 (
            .O(N__14351),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052));
    CascadeMux I__3105 (
            .O(N__14344),
            .I(N__14341));
    InMux I__3104 (
            .O(N__14341),
            .I(N__14338));
    LocalMux I__3103 (
            .O(N__14338),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i));
    InMux I__3102 (
            .O(N__14335),
            .I(N__14332));
    LocalMux I__3101 (
            .O(N__14332),
            .I(N__14329));
    Glb2LocalMux I__3100 (
            .O(N__14329),
            .I(N__14314));
    ClkMux I__3099 (
            .O(N__14328),
            .I(N__14314));
    ClkMux I__3098 (
            .O(N__14327),
            .I(N__14314));
    ClkMux I__3097 (
            .O(N__14326),
            .I(N__14314));
    ClkMux I__3096 (
            .O(N__14325),
            .I(N__14314));
    GlobalMux I__3095 (
            .O(N__14314),
            .I(N__14311));
    gio2CtrlBuf I__3094 (
            .O(N__14311),
            .I(Clock12MHz_c_g));
    IoInMux I__3093 (
            .O(N__14308),
            .I(N__14303));
    IoInMux I__3092 (
            .O(N__14307),
            .I(N__14300));
    IoInMux I__3091 (
            .O(N__14306),
            .I(N__14297));
    LocalMux I__3090 (
            .O(N__14303),
            .I(N__14292));
    LocalMux I__3089 (
            .O(N__14300),
            .I(N__14292));
    LocalMux I__3088 (
            .O(N__14297),
            .I(N__14289));
    Span12Mux_s11_v I__3087 (
            .O(N__14292),
            .I(N__14286));
    Span12Mux_s10_h I__3086 (
            .O(N__14289),
            .I(N__14283));
    Odrv12 I__3085 (
            .O(N__14286),
            .I(GB_BUFFER_Clock12MHz_c_g_THRU_CO));
    Odrv12 I__3084 (
            .O(N__14283),
            .I(GB_BUFFER_Clock12MHz_c_g_THRU_CO));
    InMux I__3083 (
            .O(N__14278),
            .I(N__14275));
    LocalMux I__3082 (
            .O(N__14275),
            .I(N__14272));
    Odrv4 I__3081 (
            .O(N__14272),
            .I(N_1557_0));
    InMux I__3080 (
            .O(N__14269),
            .I(N__14266));
    LocalMux I__3079 (
            .O(N__14266),
            .I(N__14263));
    Odrv12 I__3078 (
            .O(N__14263),
            .I(N_41_0_0_0));
    CascadeMux I__3077 (
            .O(N__14260),
            .I(N__14257));
    InMux I__3076 (
            .O(N__14257),
            .I(N__14250));
    CascadeMux I__3075 (
            .O(N__14256),
            .I(N__14247));
    InMux I__3074 (
            .O(N__14255),
            .I(N__14241));
    CascadeMux I__3073 (
            .O(N__14254),
            .I(N__14234));
    CascadeMux I__3072 (
            .O(N__14253),
            .I(N__14231));
    LocalMux I__3071 (
            .O(N__14250),
            .I(N__14228));
    InMux I__3070 (
            .O(N__14247),
            .I(N__14225));
    CascadeMux I__3069 (
            .O(N__14246),
            .I(N__14222));
    CascadeMux I__3068 (
            .O(N__14245),
            .I(N__14218));
    CascadeMux I__3067 (
            .O(N__14244),
            .I(N__14214));
    LocalMux I__3066 (
            .O(N__14241),
            .I(N__14211));
    InMux I__3065 (
            .O(N__14240),
            .I(N__14206));
    InMux I__3064 (
            .O(N__14239),
            .I(N__14206));
    InMux I__3063 (
            .O(N__14238),
            .I(N__14203));
    InMux I__3062 (
            .O(N__14237),
            .I(N__14196));
    InMux I__3061 (
            .O(N__14234),
            .I(N__14196));
    InMux I__3060 (
            .O(N__14231),
            .I(N__14196));
    Span4Mux_v I__3059 (
            .O(N__14228),
            .I(N__14191));
    LocalMux I__3058 (
            .O(N__14225),
            .I(N__14191));
    InMux I__3057 (
            .O(N__14222),
            .I(N__14184));
    InMux I__3056 (
            .O(N__14221),
            .I(N__14184));
    InMux I__3055 (
            .O(N__14218),
            .I(N__14184));
    InMux I__3054 (
            .O(N__14217),
            .I(N__14179));
    InMux I__3053 (
            .O(N__14214),
            .I(N__14179));
    Odrv4 I__3052 (
            .O(N__14211),
            .I(N_563));
    LocalMux I__3051 (
            .O(N__14206),
            .I(N_563));
    LocalMux I__3050 (
            .O(N__14203),
            .I(N_563));
    LocalMux I__3049 (
            .O(N__14196),
            .I(N_563));
    Odrv4 I__3048 (
            .O(N__14191),
            .I(N_563));
    LocalMux I__3047 (
            .O(N__14184),
            .I(N_563));
    LocalMux I__3046 (
            .O(N__14179),
            .I(N_563));
    CascadeMux I__3045 (
            .O(N__14164),
            .I(un116_pixel_5_bmZ0Z_5_cascade_));
    InMux I__3044 (
            .O(N__14161),
            .I(N__14158));
    LocalMux I__3043 (
            .O(N__14158),
            .I(N__14155));
    Span4Mux_h I__3042 (
            .O(N__14155),
            .I(N__14152));
    Odrv4 I__3041 (
            .O(N__14152),
            .I(un116_pixel_6_ns_1_5));
    InMux I__3040 (
            .O(N__14149),
            .I(N__14146));
    LocalMux I__3039 (
            .O(N__14146),
            .I(if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx));
    CascadeMux I__3038 (
            .O(N__14143),
            .I(N__14140));
    InMux I__3037 (
            .O(N__14140),
            .I(N__14137));
    LocalMux I__3036 (
            .O(N__14137),
            .I(N_858_i));
    CascadeMux I__3035 (
            .O(N__14134),
            .I(N__14131));
    InMux I__3034 (
            .O(N__14131),
            .I(N__14128));
    LocalMux I__3033 (
            .O(N__14128),
            .I(N__14125));
    Odrv4 I__3032 (
            .O(N__14125),
            .I(column_1_if_generate_plus_mult1_un47_sum1_3));
    InMux I__3031 (
            .O(N__14122),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_2));
    CascadeMux I__3030 (
            .O(N__14119),
            .I(N__14116));
    InMux I__3029 (
            .O(N__14116),
            .I(N__14113));
    LocalMux I__3028 (
            .O(N__14113),
            .I(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx));
    InMux I__3027 (
            .O(N__14110),
            .I(N__14107));
    LocalMux I__3026 (
            .O(N__14107),
            .I(column_1_if_generate_plus_mult1_un47_sum1_4));
    InMux I__3025 (
            .O(N__14104),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_3));
    InMux I__3024 (
            .O(N__14101),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_4));
    CascadeMux I__3023 (
            .O(N__14098),
            .I(N__14094));
    CascadeMux I__3022 (
            .O(N__14097),
            .I(N__14090));
    InMux I__3021 (
            .O(N__14094),
            .I(N__14086));
    InMux I__3020 (
            .O(N__14093),
            .I(N__14079));
    InMux I__3019 (
            .O(N__14090),
            .I(N__14079));
    InMux I__3018 (
            .O(N__14089),
            .I(N__14079));
    LocalMux I__3017 (
            .O(N__14086),
            .I(column_1_if_generate_plus_mult1_un47_sum1_5));
    LocalMux I__3016 (
            .O(N__14079),
            .I(column_1_if_generate_plus_mult1_un47_sum1_5));
    CascadeMux I__3015 (
            .O(N__14074),
            .I(N__14070));
    CascadeMux I__3014 (
            .O(N__14073),
            .I(N__14067));
    InMux I__3013 (
            .O(N__14070),
            .I(N__14062));
    InMux I__3012 (
            .O(N__14067),
            .I(N__14062));
    LocalMux I__3011 (
            .O(N__14062),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8));
    InMux I__3010 (
            .O(N__14059),
            .I(N__14054));
    InMux I__3009 (
            .O(N__14058),
            .I(N__14049));
    InMux I__3008 (
            .O(N__14057),
            .I(N__14049));
    LocalMux I__3007 (
            .O(N__14054),
            .I(N__14043));
    LocalMux I__3006 (
            .O(N__14049),
            .I(N__14043));
    InMux I__3005 (
            .O(N__14048),
            .I(N__14040));
    Span4Mux_v I__3004 (
            .O(N__14043),
            .I(N__14033));
    LocalMux I__3003 (
            .O(N__14040),
            .I(N__14033));
    InMux I__3002 (
            .O(N__14039),
            .I(N__14025));
    InMux I__3001 (
            .O(N__14038),
            .I(N__14025));
    Span4Mux_h I__3000 (
            .O(N__14033),
            .I(N__14022));
    InMux I__2999 (
            .O(N__14032),
            .I(N__14017));
    InMux I__2998 (
            .O(N__14031),
            .I(N__14017));
    InMux I__2997 (
            .O(N__14030),
            .I(N__14014));
    LocalMux I__2996 (
            .O(N__14025),
            .I(charx_if_generate_plus_mult1_un33_sum));
    Odrv4 I__2995 (
            .O(N__14022),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__2994 (
            .O(N__14017),
            .I(charx_if_generate_plus_mult1_un33_sum));
    LocalMux I__2993 (
            .O(N__14014),
            .I(charx_if_generate_plus_mult1_un33_sum));
    CascadeMux I__2992 (
            .O(N__14005),
            .I(N__14000));
    InMux I__2991 (
            .O(N__14004),
            .I(N__13995));
    InMux I__2990 (
            .O(N__14003),
            .I(N__13995));
    InMux I__2989 (
            .O(N__14000),
            .I(N__13992));
    LocalMux I__2988 (
            .O(N__13995),
            .I(N__13989));
    LocalMux I__2987 (
            .O(N__13992),
            .I(N_66));
    Odrv4 I__2986 (
            .O(N__13989),
            .I(N_66));
    CascadeMux I__2985 (
            .O(N__13984),
            .I(N__13981));
    InMux I__2984 (
            .O(N__13981),
            .I(N__13978));
    LocalMux I__2983 (
            .O(N__13978),
            .I(N__13975));
    Odrv4 I__2982 (
            .O(N__13975),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5LZ0));
    InMux I__2981 (
            .O(N__13972),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__2980 (
            .O(N__13969),
            .I(N__13966));
    LocalMux I__2979 (
            .O(N__13966),
            .I(N__13963));
    Odrv4 I__2978 (
            .O(N__13963),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7JZ0Z31));
    InMux I__2977 (
            .O(N__13960),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__2976 (
            .O(N__13957),
            .I(N__13954));
    LocalMux I__2975 (
            .O(N__13954),
            .I(N__13951));
    Odrv12 I__2974 (
            .O(N__13951),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUHZ0Z2));
    InMux I__2973 (
            .O(N__13948),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__2972 (
            .O(N__13945),
            .I(N__13942));
    InMux I__2971 (
            .O(N__13942),
            .I(N__13939));
    LocalMux I__2970 (
            .O(N__13939),
            .I(N__13936));
    Odrv12 I__2969 (
            .O(N__13936),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIVZ0Z6153));
    InMux I__2968 (
            .O(N__13933),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__2967 (
            .O(N__13930),
            .I(N__13927));
    LocalMux I__2966 (
            .O(N__13927),
            .I(N__13924));
    Odrv12 I__2965 (
            .O(N__13924),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__2964 (
            .O(N__13921),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__2963 (
            .O(N__13918),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7));
    CascadeMux I__2962 (
            .O(N__13915),
            .I(N__13912));
    InMux I__2961 (
            .O(N__13912),
            .I(N__13905));
    InMux I__2960 (
            .O(N__13911),
            .I(N__13905));
    InMux I__2959 (
            .O(N__13910),
            .I(N__13902));
    LocalMux I__2958 (
            .O(N__13905),
            .I(N__13899));
    LocalMux I__2957 (
            .O(N__13902),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3));
    Odrv12 I__2956 (
            .O(N__13899),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3));
    InMux I__2955 (
            .O(N__13894),
            .I(N__13891));
    LocalMux I__2954 (
            .O(N__13891),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i));
    InMux I__2953 (
            .O(N__13888),
            .I(N__13882));
    InMux I__2952 (
            .O(N__13887),
            .I(N__13877));
    InMux I__2951 (
            .O(N__13886),
            .I(N__13877));
    InMux I__2950 (
            .O(N__13885),
            .I(N__13873));
    LocalMux I__2949 (
            .O(N__13882),
            .I(N__13869));
    LocalMux I__2948 (
            .O(N__13877),
            .I(N__13865));
    InMux I__2947 (
            .O(N__13876),
            .I(N__13862));
    LocalMux I__2946 (
            .O(N__13873),
            .I(N__13859));
    InMux I__2945 (
            .O(N__13872),
            .I(N__13855));
    Span4Mux_h I__2944 (
            .O(N__13869),
            .I(N__13852));
    InMux I__2943 (
            .O(N__13868),
            .I(N__13849));
    Span4Mux_h I__2942 (
            .O(N__13865),
            .I(N__13842));
    LocalMux I__2941 (
            .O(N__13862),
            .I(N__13842));
    Span4Mux_h I__2940 (
            .O(N__13859),
            .I(N__13842));
    InMux I__2939 (
            .O(N__13858),
            .I(N__13839));
    LocalMux I__2938 (
            .O(N__13855),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2937 (
            .O(N__13852),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__2936 (
            .O(N__13849),
            .I(charx_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2935 (
            .O(N__13842),
            .I(charx_if_generate_plus_mult1_un40_sum));
    LocalMux I__2934 (
            .O(N__13839),
            .I(charx_if_generate_plus_mult1_un40_sum));
    CascadeMux I__2933 (
            .O(N__13828),
            .I(N__13825));
    InMux I__2932 (
            .O(N__13825),
            .I(N__13822));
    LocalMux I__2931 (
            .O(N__13822),
            .I(un5_visiblex_i_0_25));
    CascadeMux I__2930 (
            .O(N__13819),
            .I(N__13816));
    InMux I__2929 (
            .O(N__13816),
            .I(N__13813));
    LocalMux I__2928 (
            .O(N__13813),
            .I(column_1_if_generate_plus_mult1_un47_sum1_2));
    InMux I__2927 (
            .O(N__13810),
            .I(column_1_if_generate_plus_mult1_un47_sum_1_cry_1));
    CascadeMux I__2926 (
            .O(N__13807),
            .I(N__13804));
    InMux I__2925 (
            .O(N__13804),
            .I(N__13801));
    LocalMux I__2924 (
            .O(N__13801),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0));
    InMux I__2923 (
            .O(N__13798),
            .I(N__13795));
    LocalMux I__2922 (
            .O(N__13795),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8TZ0Z77));
    InMux I__2921 (
            .O(N__13792),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1));
    CascadeMux I__2920 (
            .O(N__13789),
            .I(N__13786));
    InMux I__2919 (
            .O(N__13786),
            .I(N__13783));
    LocalMux I__2918 (
            .O(N__13783),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0));
    InMux I__2917 (
            .O(N__13780),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2));
    CascadeMux I__2916 (
            .O(N__13777),
            .I(N__13773));
    InMux I__2915 (
            .O(N__13776),
            .I(N__13770));
    InMux I__2914 (
            .O(N__13773),
            .I(N__13767));
    LocalMux I__2913 (
            .O(N__13770),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    LocalMux I__2912 (
            .O(N__13767),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf));
    InMux I__2911 (
            .O(N__13762),
            .I(N__13759));
    LocalMux I__2910 (
            .O(N__13759),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO));
    InMux I__2909 (
            .O(N__13756),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3));
    InMux I__2908 (
            .O(N__13753),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4));
    InMux I__2907 (
            .O(N__13750),
            .I(N__13741));
    InMux I__2906 (
            .O(N__13749),
            .I(N__13741));
    InMux I__2905 (
            .O(N__13748),
            .I(N__13741));
    LocalMux I__2904 (
            .O(N__13741),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO));
    CascadeMux I__2903 (
            .O(N__13738),
            .I(N__13735));
    InMux I__2902 (
            .O(N__13735),
            .I(N__13732));
    LocalMux I__2901 (
            .O(N__13732),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77Z0Z_0));
    CascadeMux I__2900 (
            .O(N__13729),
            .I(N__13726));
    InMux I__2899 (
            .O(N__13726),
            .I(N__13723));
    LocalMux I__2898 (
            .O(N__13723),
            .I(charx_i_23));
    CascadeMux I__2897 (
            .O(N__13720),
            .I(N__13716));
    InMux I__2896 (
            .O(N__13719),
            .I(N__13710));
    InMux I__2895 (
            .O(N__13716),
            .I(N__13705));
    InMux I__2894 (
            .O(N__13715),
            .I(N__13705));
    InMux I__2893 (
            .O(N__13714),
            .I(N__13702));
    InMux I__2892 (
            .O(N__13713),
            .I(N__13699));
    LocalMux I__2891 (
            .O(N__13710),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1));
    LocalMux I__2890 (
            .O(N__13705),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1));
    LocalMux I__2889 (
            .O(N__13702),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1));
    LocalMux I__2888 (
            .O(N__13699),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1));
    CascadeMux I__2887 (
            .O(N__13690),
            .I(N__13685));
    CascadeMux I__2886 (
            .O(N__13689),
            .I(N__13682));
    CascadeMux I__2885 (
            .O(N__13688),
            .I(N__13679));
    InMux I__2884 (
            .O(N__13685),
            .I(N__13676));
    InMux I__2883 (
            .O(N__13682),
            .I(N__13673));
    InMux I__2882 (
            .O(N__13679),
            .I(N__13670));
    LocalMux I__2881 (
            .O(N__13676),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2));
    LocalMux I__2880 (
            .O(N__13673),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2));
    LocalMux I__2879 (
            .O(N__13670),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2));
    InMux I__2878 (
            .O(N__13663),
            .I(N__13660));
    LocalMux I__2877 (
            .O(N__13660),
            .I(N__13653));
    InMux I__2876 (
            .O(N__13659),
            .I(N__13650));
    InMux I__2875 (
            .O(N__13658),
            .I(N__13645));
    InMux I__2874 (
            .O(N__13657),
            .I(N__13645));
    InMux I__2873 (
            .O(N__13656),
            .I(N__13642));
    Odrv4 I__2872 (
            .O(N__13653),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843));
    LocalMux I__2871 (
            .O(N__13650),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843));
    LocalMux I__2870 (
            .O(N__13645),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843));
    LocalMux I__2869 (
            .O(N__13642),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843));
    CascadeMux I__2868 (
            .O(N__13633),
            .I(N__13630));
    InMux I__2867 (
            .O(N__13630),
            .I(N__13627));
    LocalMux I__2866 (
            .O(N__13627),
            .I(charx_i_24));
    InMux I__2865 (
            .O(N__13624),
            .I(N__13621));
    LocalMux I__2864 (
            .O(N__13621),
            .I(un116_pixel_2_bm_0));
    InMux I__2863 (
            .O(N__13618),
            .I(N__13615));
    LocalMux I__2862 (
            .O(N__13615),
            .I(un114_pixel_1_0_3__un116_pixel_5_ns_1_0Z0Z_0));
    CascadeMux I__2861 (
            .O(N__13612),
            .I(N__13608));
    InMux I__2860 (
            .O(N__13611),
            .I(N__13604));
    InMux I__2859 (
            .O(N__13608),
            .I(N__13600));
    InMux I__2858 (
            .O(N__13607),
            .I(N__13596));
    LocalMux I__2857 (
            .O(N__13604),
            .I(N__13593));
    InMux I__2856 (
            .O(N__13603),
            .I(N__13590));
    LocalMux I__2855 (
            .O(N__13600),
            .I(N__13587));
    InMux I__2854 (
            .O(N__13599),
            .I(N__13584));
    LocalMux I__2853 (
            .O(N__13596),
            .I(N__13581));
    Span4Mux_v I__2852 (
            .O(N__13593),
            .I(N__13578));
    LocalMux I__2851 (
            .O(N__13590),
            .I(N__13575));
    Span4Mux_h I__2850 (
            .O(N__13587),
            .I(N__13572));
    LocalMux I__2849 (
            .O(N__13584),
            .I(N__13569));
    Span4Mux_v I__2848 (
            .O(N__13581),
            .I(N__13564));
    Span4Mux_s3_h I__2847 (
            .O(N__13578),
            .I(N__13564));
    Span4Mux_s3_v I__2846 (
            .O(N__13575),
            .I(N__13561));
    Odrv4 I__2845 (
            .O(N__13572),
            .I(chessboardpixel_un152_pixel_24));
    Odrv4 I__2844 (
            .O(N__13569),
            .I(chessboardpixel_un152_pixel_24));
    Odrv4 I__2843 (
            .O(N__13564),
            .I(chessboardpixel_un152_pixel_24));
    Odrv4 I__2842 (
            .O(N__13561),
            .I(chessboardpixel_un152_pixel_24));
    InMux I__2841 (
            .O(N__13552),
            .I(N__13549));
    LocalMux I__2840 (
            .O(N__13549),
            .I(N__13546));
    Odrv4 I__2839 (
            .O(N__13546),
            .I(un114_pixel_1_0_3__un116_pixel_6_1_1Z0Z_1));
    InMux I__2838 (
            .O(N__13543),
            .I(N__13537));
    InMux I__2837 (
            .O(N__13542),
            .I(N__13533));
    InMux I__2836 (
            .O(N__13541),
            .I(N__13528));
    InMux I__2835 (
            .O(N__13540),
            .I(N__13528));
    LocalMux I__2834 (
            .O(N__13537),
            .I(N__13525));
    InMux I__2833 (
            .O(N__13536),
            .I(N__13522));
    LocalMux I__2832 (
            .O(N__13533),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__2831 (
            .O(N__13528),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    Odrv4 I__2830 (
            .O(N__13525),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    LocalMux I__2829 (
            .O(N__13522),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1));
    CascadeMux I__2828 (
            .O(N__13513),
            .I(N__13510));
    InMux I__2827 (
            .O(N__13510),
            .I(N__13506));
    InMux I__2826 (
            .O(N__13509),
            .I(N__13503));
    LocalMux I__2825 (
            .O(N__13506),
            .I(N__13500));
    LocalMux I__2824 (
            .O(N__13503),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4));
    Odrv4 I__2823 (
            .O(N__13500),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4));
    InMux I__2822 (
            .O(N__13495),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1));
    InMux I__2821 (
            .O(N__13492),
            .I(N__13489));
    LocalMux I__2820 (
            .O(N__13489),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3EZ0Z987));
    InMux I__2819 (
            .O(N__13486),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2));
    CascadeMux I__2818 (
            .O(N__13483),
            .I(N__13479));
    CascadeMux I__2817 (
            .O(N__13482),
            .I(N__13476));
    InMux I__2816 (
            .O(N__13479),
            .I(N__13471));
    InMux I__2815 (
            .O(N__13476),
            .I(N__13471));
    LocalMux I__2814 (
            .O(N__13471),
            .I(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803));
    InMux I__2813 (
            .O(N__13468),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4));
    CascadeMux I__2812 (
            .O(N__13465),
            .I(N__13461));
    InMux I__2811 (
            .O(N__13464),
            .I(N__13455));
    InMux I__2810 (
            .O(N__13461),
            .I(N__13452));
    InMux I__2809 (
            .O(N__13460),
            .I(N__13449));
    InMux I__2808 (
            .O(N__13459),
            .I(N__13444));
    InMux I__2807 (
            .O(N__13458),
            .I(N__13444));
    LocalMux I__2806 (
            .O(N__13455),
            .I(N__13441));
    LocalMux I__2805 (
            .O(N__13452),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987));
    LocalMux I__2804 (
            .O(N__13449),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987));
    LocalMux I__2803 (
            .O(N__13444),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987));
    Odrv4 I__2802 (
            .O(N__13441),
            .I(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987));
    InMux I__2801 (
            .O(N__13432),
            .I(N__13429));
    LocalMux I__2800 (
            .O(N__13429),
            .I(un116_pixel_4_am_1));
    CascadeMux I__2799 (
            .O(N__13426),
            .I(N__13419));
    InMux I__2798 (
            .O(N__13425),
            .I(N__13414));
    InMux I__2797 (
            .O(N__13424),
            .I(N__13409));
    InMux I__2796 (
            .O(N__13423),
            .I(N__13409));
    InMux I__2795 (
            .O(N__13422),
            .I(N__13406));
    InMux I__2794 (
            .O(N__13419),
            .I(N__13403));
    InMux I__2793 (
            .O(N__13418),
            .I(N__13400));
    InMux I__2792 (
            .O(N__13417),
            .I(N__13397));
    LocalMux I__2791 (
            .O(N__13414),
            .I(N__13394));
    LocalMux I__2790 (
            .O(N__13409),
            .I(N_36));
    LocalMux I__2789 (
            .O(N__13406),
            .I(N_36));
    LocalMux I__2788 (
            .O(N__13403),
            .I(N_36));
    LocalMux I__2787 (
            .O(N__13400),
            .I(N_36));
    LocalMux I__2786 (
            .O(N__13397),
            .I(N_36));
    Odrv4 I__2785 (
            .O(N__13394),
            .I(N_36));
    InMux I__2784 (
            .O(N__13381),
            .I(N__13378));
    LocalMux I__2783 (
            .O(N__13378),
            .I(un116_pixel_5_amZ0Z_5));
    InMux I__2782 (
            .O(N__13375),
            .I(N__13372));
    LocalMux I__2781 (
            .O(N__13372),
            .I(un116_pixel_2_amZ0Z_5));
    InMux I__2780 (
            .O(N__13369),
            .I(N__13366));
    LocalMux I__2779 (
            .O(N__13366),
            .I(N_385));
    InMux I__2778 (
            .O(N__13363),
            .I(N__13359));
    InMux I__2777 (
            .O(N__13362),
            .I(N__13356));
    LocalMux I__2776 (
            .O(N__13359),
            .I(N_325));
    LocalMux I__2775 (
            .O(N__13356),
            .I(N_325));
    InMux I__2774 (
            .O(N__13351),
            .I(N__13348));
    LocalMux I__2773 (
            .O(N__13348),
            .I(un116_pixel_2_bmZ0Z_1));
    InMux I__2772 (
            .O(N__13345),
            .I(N__13342));
    LocalMux I__2771 (
            .O(N__13342),
            .I(un114_pixel_1_0_3__un116_pixel_6_1Z0Z_1));
    InMux I__2770 (
            .O(N__13339),
            .I(N__13336));
    LocalMux I__2769 (
            .O(N__13336),
            .I(N__13331));
    InMux I__2768 (
            .O(N__13335),
            .I(N__13328));
    InMux I__2767 (
            .O(N__13334),
            .I(N__13325));
    Odrv4 I__2766 (
            .O(N__13331),
            .I(un116_pixel_1_4));
    LocalMux I__2765 (
            .O(N__13328),
            .I(un116_pixel_1_4));
    LocalMux I__2764 (
            .O(N__13325),
            .I(un116_pixel_1_4));
    InMux I__2763 (
            .O(N__13318),
            .I(N__13314));
    InMux I__2762 (
            .O(N__13317),
            .I(N__13311));
    LocalMux I__2761 (
            .O(N__13314),
            .I(N_374_0));
    LocalMux I__2760 (
            .O(N__13311),
            .I(N_374_0));
    CascadeMux I__2759 (
            .O(N__13306),
            .I(N__13296));
    InMux I__2758 (
            .O(N__13305),
            .I(N__13285));
    InMux I__2757 (
            .O(N__13304),
            .I(N__13285));
    InMux I__2756 (
            .O(N__13303),
            .I(N__13285));
    InMux I__2755 (
            .O(N__13302),
            .I(N__13282));
    InMux I__2754 (
            .O(N__13301),
            .I(N__13275));
    InMux I__2753 (
            .O(N__13300),
            .I(N__13275));
    InMux I__2752 (
            .O(N__13299),
            .I(N__13275));
    InMux I__2751 (
            .O(N__13296),
            .I(N__13270));
    InMux I__2750 (
            .O(N__13295),
            .I(N__13270));
    InMux I__2749 (
            .O(N__13294),
            .I(N__13267));
    InMux I__2748 (
            .O(N__13293),
            .I(N__13262));
    InMux I__2747 (
            .O(N__13292),
            .I(N__13262));
    LocalMux I__2746 (
            .O(N__13285),
            .I(font_un3_pixel_29));
    LocalMux I__2745 (
            .O(N__13282),
            .I(font_un3_pixel_29));
    LocalMux I__2744 (
            .O(N__13275),
            .I(font_un3_pixel_29));
    LocalMux I__2743 (
            .O(N__13270),
            .I(font_un3_pixel_29));
    LocalMux I__2742 (
            .O(N__13267),
            .I(font_un3_pixel_29));
    LocalMux I__2741 (
            .O(N__13262),
            .I(font_un3_pixel_29));
    CascadeMux I__2740 (
            .O(N__13249),
            .I(un116_pixel_7_x0_0_cascade_));
    InMux I__2739 (
            .O(N__13246),
            .I(N__13243));
    LocalMux I__2738 (
            .O(N__13243),
            .I(un116_pixel_7_x1_0));
    InMux I__2737 (
            .O(N__13240),
            .I(N__13237));
    LocalMux I__2736 (
            .O(N__13237),
            .I(un116_pixel_7_ns_0));
    InMux I__2735 (
            .O(N__13234),
            .I(N__13231));
    LocalMux I__2734 (
            .O(N__13231),
            .I(column_0111_0));
    InMux I__2733 (
            .O(N__13228),
            .I(N__13225));
    LocalMux I__2732 (
            .O(N__13225),
            .I(un116_pixel_3_ns_1_0_3));
    InMux I__2731 (
            .O(N__13222),
            .I(N__13219));
    LocalMux I__2730 (
            .O(N__13219),
            .I(un114_pixel_1_0_3__g1Z0Z_4));
    CascadeMux I__2729 (
            .O(N__13216),
            .I(N_1583_0_cascade_));
    InMux I__2728 (
            .O(N__13213),
            .I(N__13210));
    LocalMux I__2727 (
            .O(N__13210),
            .I(N_26_0_0));
    CascadeMux I__2726 (
            .O(N__13207),
            .I(un116_pixel_2_amZ0Z_1_cascade_));
    InMux I__2725 (
            .O(N__13204),
            .I(N__13201));
    LocalMux I__2724 (
            .O(N__13201),
            .I(un116_pixel_6_1));
    CascadeMux I__2723 (
            .O(N__13198),
            .I(column_0001_0_cascade_));
    InMux I__2722 (
            .O(N__13195),
            .I(N__13192));
    LocalMux I__2721 (
            .O(N__13192),
            .I(beamY_RNILBST4T2Z0Z_1));
    CascadeMux I__2720 (
            .O(N__13189),
            .I(beamY_RNIT81CMJ2Z0Z_1_cascade_));
    InMux I__2719 (
            .O(N__13186),
            .I(N__13183));
    LocalMux I__2718 (
            .O(N__13183),
            .I(N__13180));
    Odrv4 I__2717 (
            .O(N__13180),
            .I(font_un126_pixel_2_am));
    InMux I__2716 (
            .O(N__13177),
            .I(N__13174));
    LocalMux I__2715 (
            .O(N__13174),
            .I(N__13171));
    Span4Mux_h I__2714 (
            .O(N__13171),
            .I(N__13168));
    Odrv4 I__2713 (
            .O(N__13168),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5RZ0));
    InMux I__2712 (
            .O(N__13165),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_1));
    InMux I__2711 (
            .O(N__13162),
            .I(N__13158));
    InMux I__2710 (
            .O(N__13161),
            .I(N__13155));
    LocalMux I__2709 (
            .O(N__13158),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0));
    LocalMux I__2708 (
            .O(N__13155),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0));
    CascadeMux I__2707 (
            .O(N__13150),
            .I(N__13147));
    InMux I__2706 (
            .O(N__13147),
            .I(N__13144));
    LocalMux I__2705 (
            .O(N__13144),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRDZ0));
    InMux I__2704 (
            .O(N__13141),
            .I(N__13138));
    LocalMux I__2703 (
            .O(N__13138),
            .I(N__13135));
    Span4Mux_h I__2702 (
            .O(N__13135),
            .I(N__13132));
    Odrv4 I__2701 (
            .O(N__13132),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BVZ0Z81));
    InMux I__2700 (
            .O(N__13129),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__2699 (
            .O(N__13126),
            .I(N__13123));
    LocalMux I__2698 (
            .O(N__13123),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0LZ0));
    CascadeMux I__2697 (
            .O(N__13120),
            .I(N__13116));
    CascadeMux I__2696 (
            .O(N__13119),
            .I(N__13113));
    InMux I__2695 (
            .O(N__13116),
            .I(N__13108));
    InMux I__2694 (
            .O(N__13113),
            .I(N__13108));
    LocalMux I__2693 (
            .O(N__13108),
            .I(charx_if_generate_plus_mult1_un61_sum_i_5));
    InMux I__2692 (
            .O(N__13105),
            .I(N__13102));
    LocalMux I__2691 (
            .O(N__13102),
            .I(N__13099));
    Span4Mux_h I__2690 (
            .O(N__13099),
            .I(N__13096));
    Odrv4 I__2689 (
            .O(N__13096),
            .I(charx_if_generate_plus_mult1_un75_sum_axb_5));
    InMux I__2688 (
            .O(N__13093),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__2687 (
            .O(N__13090),
            .I(N__13087));
    LocalMux I__2686 (
            .O(N__13087),
            .I(charx_if_generate_plus_mult1_un68_sum_axb_5));
    InMux I__2685 (
            .O(N__13084),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__2684 (
            .O(N__13081),
            .I(N__13078));
    InMux I__2683 (
            .O(N__13078),
            .I(N__13071));
    InMux I__2682 (
            .O(N__13077),
            .I(N__13071));
    InMux I__2681 (
            .O(N__13076),
            .I(N__13067));
    LocalMux I__2680 (
            .O(N__13071),
            .I(N__13064));
    InMux I__2679 (
            .O(N__13070),
            .I(N__13061));
    LocalMux I__2678 (
            .O(N__13067),
            .I(N__13056));
    Span4Mux_h I__2677 (
            .O(N__13064),
            .I(N__13056));
    LocalMux I__2676 (
            .O(N__13061),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1));
    Odrv4 I__2675 (
            .O(N__13056),
            .I(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1));
    InMux I__2674 (
            .O(N__13051),
            .I(N__13048));
    LocalMux I__2673 (
            .O(N__13048),
            .I(charx_if_generate_plus_mult1_un61_sum_i));
    InMux I__2672 (
            .O(N__13045),
            .I(N__13042));
    LocalMux I__2671 (
            .O(N__13042),
            .I(N_41_0));
    CascadeMux I__2670 (
            .O(N__13039),
            .I(column_1_if_generate_plus_mult1_un54_sum_axb_2_sxZ0_cascade_));
    CascadeMux I__2669 (
            .O(N__13036),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2_cascade_));
    InMux I__2668 (
            .O(N__13033),
            .I(N__13030));
    LocalMux I__2667 (
            .O(N__13030),
            .I(if_generate_plus_mult1_un54_sum_axb_2_l_fx));
    InMux I__2666 (
            .O(N__13027),
            .I(N__13024));
    LocalMux I__2665 (
            .O(N__13024),
            .I(column_1_if_generate_plus_mult1_un47_sum0_4));
    CascadeMux I__2664 (
            .O(N__13021),
            .I(if_generate_plus_mult1_un47_sum_m_5_cascade_));
    InMux I__2663 (
            .O(N__13018),
            .I(N__13015));
    LocalMux I__2662 (
            .O(N__13015),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5));
    InMux I__2661 (
            .O(N__13012),
            .I(N__13009));
    LocalMux I__2660 (
            .O(N__13009),
            .I(column_1_if_generate_plus_mult1_un47_sum0_2));
    InMux I__2659 (
            .O(N__13006),
            .I(N__13001));
    InMux I__2658 (
            .O(N__13005),
            .I(N__12996));
    InMux I__2657 (
            .O(N__13004),
            .I(N__12996));
    LocalMux I__2656 (
            .O(N__13001),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    LocalMux I__2655 (
            .O(N__12996),
            .I(if_generate_plus_mult1_un47_sum_m_5));
    CascadeMux I__2654 (
            .O(N__12991),
            .I(N__12988));
    InMux I__2653 (
            .O(N__12988),
            .I(N__12985));
    LocalMux I__2652 (
            .O(N__12985),
            .I(if_generate_plus_mult1_un54_sum_axb_3_l_fx));
    InMux I__2651 (
            .O(N__12982),
            .I(N__12976));
    InMux I__2650 (
            .O(N__12981),
            .I(N__12969));
    InMux I__2649 (
            .O(N__12980),
            .I(N__12969));
    InMux I__2648 (
            .O(N__12979),
            .I(N__12969));
    LocalMux I__2647 (
            .O(N__12976),
            .I(column_1_if_generate_plus_mult1_un47_sum0_5));
    LocalMux I__2646 (
            .O(N__12969),
            .I(column_1_if_generate_plus_mult1_un47_sum0_5));
    CascadeMux I__2645 (
            .O(N__12964),
            .I(N__12960));
    CascadeMux I__2644 (
            .O(N__12963),
            .I(N__12957));
    InMux I__2643 (
            .O(N__12960),
            .I(N__12950));
    InMux I__2642 (
            .O(N__12957),
            .I(N__12950));
    InMux I__2641 (
            .O(N__12956),
            .I(N__12947));
    InMux I__2640 (
            .O(N__12955),
            .I(N__12944));
    LocalMux I__2639 (
            .O(N__12950),
            .I(N_584_i));
    LocalMux I__2638 (
            .O(N__12947),
            .I(N_584_i));
    LocalMux I__2637 (
            .O(N__12944),
            .I(N_584_i));
    InMux I__2636 (
            .O(N__12937),
            .I(N__12931));
    InMux I__2635 (
            .O(N__12936),
            .I(N__12928));
    CascadeMux I__2634 (
            .O(N__12935),
            .I(N__12925));
    CascadeMux I__2633 (
            .O(N__12934),
            .I(N__12920));
    LocalMux I__2632 (
            .O(N__12931),
            .I(N__12915));
    LocalMux I__2631 (
            .O(N__12928),
            .I(N__12912));
    InMux I__2630 (
            .O(N__12925),
            .I(N__12907));
    InMux I__2629 (
            .O(N__12924),
            .I(N__12907));
    InMux I__2628 (
            .O(N__12923),
            .I(N__12902));
    InMux I__2627 (
            .O(N__12920),
            .I(N__12902));
    InMux I__2626 (
            .O(N__12919),
            .I(N__12897));
    InMux I__2625 (
            .O(N__12918),
            .I(N__12897));
    Span4Mux_h I__2624 (
            .O(N__12915),
            .I(N__12885));
    Span4Mux_v I__2623 (
            .O(N__12912),
            .I(N__12885));
    LocalMux I__2622 (
            .O(N__12907),
            .I(N__12885));
    LocalMux I__2621 (
            .O(N__12902),
            .I(N__12885));
    LocalMux I__2620 (
            .O(N__12897),
            .I(N__12885));
    InMux I__2619 (
            .O(N__12896),
            .I(N__12882));
    Odrv4 I__2618 (
            .O(N__12885),
            .I(N_37_i));
    LocalMux I__2617 (
            .O(N__12882),
            .I(N_37_i));
    InMux I__2616 (
            .O(N__12877),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__2615 (
            .O(N__12874),
            .I(N__12871));
    InMux I__2614 (
            .O(N__12871),
            .I(N__12868));
    LocalMux I__2613 (
            .O(N__12868),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_invZ0));
    InMux I__2612 (
            .O(N__12865),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__2611 (
            .O(N__12862),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843_cascade_));
    InMux I__2610 (
            .O(N__12859),
            .I(N__12856));
    LocalMux I__2609 (
            .O(N__12856),
            .I(charx_if_generate_plus_mult1_un68_sum_i));
    CascadeMux I__2608 (
            .O(N__12853),
            .I(N__12850));
    InMux I__2607 (
            .O(N__12850),
            .I(N__12847));
    LocalMux I__2606 (
            .O(N__12847),
            .I(N__12844));
    Odrv4 I__2605 (
            .O(N__12844),
            .I(un114_pixel_1_0_3__un4_row_8Z0Z_0));
    CascadeMux I__2604 (
            .O(N__12841),
            .I(N__12838));
    InMux I__2603 (
            .O(N__12838),
            .I(N__12835));
    LocalMux I__2602 (
            .O(N__12835),
            .I(charx_if_generate_plus_mult1_un68_sum_i_5));
    InMux I__2601 (
            .O(N__12832),
            .I(N__12829));
    LocalMux I__2600 (
            .O(N__12829),
            .I(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx));
    InMux I__2599 (
            .O(N__12826),
            .I(N__12823));
    LocalMux I__2598 (
            .O(N__12823),
            .I(un114_pixel_1_0_3__font_un57_pixelZ0Z_0));
    InMux I__2597 (
            .O(N__12820),
            .I(N__12817));
    LocalMux I__2596 (
            .O(N__12817),
            .I(N__12813));
    InMux I__2595 (
            .O(N__12816),
            .I(N__12806));
    Span4Mux_v I__2594 (
            .O(N__12813),
            .I(N__12801));
    InMux I__2593 (
            .O(N__12812),
            .I(N__12798));
    InMux I__2592 (
            .O(N__12811),
            .I(N__12793));
    InMux I__2591 (
            .O(N__12810),
            .I(N__12793));
    CascadeMux I__2590 (
            .O(N__12809),
            .I(N__12788));
    LocalMux I__2589 (
            .O(N__12806),
            .I(N__12785));
    InMux I__2588 (
            .O(N__12805),
            .I(N__12782));
    CascadeMux I__2587 (
            .O(N__12804),
            .I(N__12779));
    Span4Mux_h I__2586 (
            .O(N__12801),
            .I(N__12772));
    LocalMux I__2585 (
            .O(N__12798),
            .I(N__12772));
    LocalMux I__2584 (
            .O(N__12793),
            .I(N__12772));
    InMux I__2583 (
            .O(N__12792),
            .I(N__12769));
    InMux I__2582 (
            .O(N__12791),
            .I(N__12766));
    InMux I__2581 (
            .O(N__12788),
            .I(N__12763));
    Span4Mux_h I__2580 (
            .O(N__12785),
            .I(N__12758));
    LocalMux I__2579 (
            .O(N__12782),
            .I(N__12758));
    InMux I__2578 (
            .O(N__12779),
            .I(N__12755));
    Span4Mux_v I__2577 (
            .O(N__12772),
            .I(N__12752));
    LocalMux I__2576 (
            .O(N__12769),
            .I(N__12749));
    LocalMux I__2575 (
            .O(N__12766),
            .I(N__12744));
    LocalMux I__2574 (
            .O(N__12763),
            .I(N__12744));
    Span4Mux_v I__2573 (
            .O(N__12758),
            .I(N__12739));
    LocalMux I__2572 (
            .O(N__12755),
            .I(N__12739));
    Odrv4 I__2571 (
            .O(N__12752),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2570 (
            .O(N__12749),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv12 I__2569 (
            .O(N__12744),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    Odrv4 I__2568 (
            .O(N__12739),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum));
    InMux I__2567 (
            .O(N__12730),
            .I(N__12727));
    LocalMux I__2566 (
            .O(N__12727),
            .I(N__12724));
    Span4Mux_h I__2565 (
            .O(N__12724),
            .I(N__12718));
    InMux I__2564 (
            .O(N__12723),
            .I(N__12715));
    InMux I__2563 (
            .O(N__12722),
            .I(N__12710));
    InMux I__2562 (
            .O(N__12721),
            .I(N__12710));
    Odrv4 I__2561 (
            .O(N__12718),
            .I(if_generate_plus_mult1_un61_sum_axbxc5));
    LocalMux I__2560 (
            .O(N__12715),
            .I(if_generate_plus_mult1_un61_sum_axbxc5));
    LocalMux I__2559 (
            .O(N__12710),
            .I(if_generate_plus_mult1_un61_sum_axbxc5));
    CascadeMux I__2558 (
            .O(N__12703),
            .I(un114_pixel_1_0_3__un4_row_8Z0Z_3_cascade_));
    InMux I__2557 (
            .O(N__12700),
            .I(N__12697));
    LocalMux I__2556 (
            .O(N__12697),
            .I(N__12694));
    Odrv4 I__2555 (
            .O(N__12694),
            .I(un114_pixel_1_0_3__un4_row_8_7Z0Z_1));
    InMux I__2554 (
            .O(N__12691),
            .I(N__12680));
    InMux I__2553 (
            .O(N__12690),
            .I(N__12680));
    InMux I__2552 (
            .O(N__12689),
            .I(N__12674));
    InMux I__2551 (
            .O(N__12688),
            .I(N__12674));
    InMux I__2550 (
            .O(N__12687),
            .I(N__12671));
    CascadeMux I__2549 (
            .O(N__12686),
            .I(N__12667));
    CascadeMux I__2548 (
            .O(N__12685),
            .I(N__12662));
    LocalMux I__2547 (
            .O(N__12680),
            .I(N__12659));
    InMux I__2546 (
            .O(N__12679),
            .I(N__12656));
    LocalMux I__2545 (
            .O(N__12674),
            .I(N__12651));
    LocalMux I__2544 (
            .O(N__12671),
            .I(N__12648));
    InMux I__2543 (
            .O(N__12670),
            .I(N__12641));
    InMux I__2542 (
            .O(N__12667),
            .I(N__12641));
    InMux I__2541 (
            .O(N__12666),
            .I(N__12641));
    InMux I__2540 (
            .O(N__12665),
            .I(N__12636));
    InMux I__2539 (
            .O(N__12662),
            .I(N__12636));
    Span4Mux_h I__2538 (
            .O(N__12659),
            .I(N__12631));
    LocalMux I__2537 (
            .O(N__12656),
            .I(N__12631));
    InMux I__2536 (
            .O(N__12655),
            .I(N__12626));
    InMux I__2535 (
            .O(N__12654),
            .I(N__12626));
    Span4Mux_v I__2534 (
            .O(N__12651),
            .I(N__12623));
    Span4Mux_h I__2533 (
            .O(N__12648),
            .I(N__12620));
    LocalMux I__2532 (
            .O(N__12641),
            .I(N__12615));
    LocalMux I__2531 (
            .O(N__12636),
            .I(N__12615));
    Span4Mux_h I__2530 (
            .O(N__12631),
            .I(N__12610));
    LocalMux I__2529 (
            .O(N__12626),
            .I(N__12610));
    Odrv4 I__2528 (
            .O(N__12623),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum));
    Odrv4 I__2527 (
            .O(N__12620),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum));
    Odrv4 I__2526 (
            .O(N__12615),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum));
    Odrv4 I__2525 (
            .O(N__12610),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum));
    InMux I__2524 (
            .O(N__12601),
            .I(N__12593));
    InMux I__2523 (
            .O(N__12600),
            .I(N__12593));
    CascadeMux I__2522 (
            .O(N__12599),
            .I(N__12588));
    CascadeMux I__2521 (
            .O(N__12598),
            .I(N__12585));
    LocalMux I__2520 (
            .O(N__12593),
            .I(N__12578));
    InMux I__2519 (
            .O(N__12592),
            .I(N__12575));
    InMux I__2518 (
            .O(N__12591),
            .I(N__12572));
    InMux I__2517 (
            .O(N__12588),
            .I(N__12567));
    InMux I__2516 (
            .O(N__12585),
            .I(N__12567));
    InMux I__2515 (
            .O(N__12584),
            .I(N__12560));
    InMux I__2514 (
            .O(N__12583),
            .I(N__12560));
    InMux I__2513 (
            .O(N__12582),
            .I(N__12560));
    InMux I__2512 (
            .O(N__12581),
            .I(N__12557));
    Span4Mux_v I__2511 (
            .O(N__12578),
            .I(N__12554));
    LocalMux I__2510 (
            .O(N__12575),
            .I(N__12551));
    LocalMux I__2509 (
            .O(N__12572),
            .I(N__12548));
    LocalMux I__2508 (
            .O(N__12567),
            .I(N__12545));
    LocalMux I__2507 (
            .O(N__12560),
            .I(N__12540));
    LocalMux I__2506 (
            .O(N__12557),
            .I(N__12540));
    Span4Mux_h I__2505 (
            .O(N__12554),
            .I(N__12533));
    Span4Mux_v I__2504 (
            .O(N__12551),
            .I(N__12533));
    Span4Mux_h I__2503 (
            .O(N__12548),
            .I(N__12530));
    Span4Mux_h I__2502 (
            .O(N__12545),
            .I(N__12525));
    Span4Mux_h I__2501 (
            .O(N__12540),
            .I(N__12525));
    InMux I__2500 (
            .O(N__12539),
            .I(N__12522));
    InMux I__2499 (
            .O(N__12538),
            .I(N__12519));
    Odrv4 I__2498 (
            .O(N__12533),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv4 I__2497 (
            .O(N__12530),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    Odrv4 I__2496 (
            .O(N__12525),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    LocalMux I__2495 (
            .O(N__12522),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    LocalMux I__2494 (
            .O(N__12519),
            .I(chary_if_generate_plus_mult1_un33_sum_axb3));
    CascadeMux I__2493 (
            .O(N__12508),
            .I(N__12504));
    InMux I__2492 (
            .O(N__12507),
            .I(N__12500));
    InMux I__2491 (
            .O(N__12504),
            .I(N__12494));
    InMux I__2490 (
            .O(N__12503),
            .I(N__12494));
    LocalMux I__2489 (
            .O(N__12500),
            .I(N__12491));
    InMux I__2488 (
            .O(N__12499),
            .I(N__12488));
    LocalMux I__2487 (
            .O(N__12494),
            .I(N__12485));
    Odrv4 I__2486 (
            .O(N__12491),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__2485 (
            .O(N__12488),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    Odrv12 I__2484 (
            .O(N__12485),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    CascadeMux I__2483 (
            .O(N__12478),
            .I(N__12475));
    InMux I__2482 (
            .O(N__12475),
            .I(N__12472));
    LocalMux I__2481 (
            .O(N__12472),
            .I(un114_pixel_1_0_3__un4_row_8Z0Z_2));
    InMux I__2480 (
            .O(N__12469),
            .I(N__12466));
    LocalMux I__2479 (
            .O(N__12466),
            .I(N__12462));
    CascadeMux I__2478 (
            .O(N__12465),
            .I(N__12459));
    Span4Mux_v I__2477 (
            .O(N__12462),
            .I(N__12456));
    InMux I__2476 (
            .O(N__12459),
            .I(N__12453));
    Odrv4 I__2475 (
            .O(N__12456),
            .I(row_1_if_generate_plus_mult1_un75_sum_cZ0Z5));
    LocalMux I__2474 (
            .O(N__12453),
            .I(row_1_if_generate_plus_mult1_un75_sum_cZ0Z5));
    InMux I__2473 (
            .O(N__12448),
            .I(N__12442));
    InMux I__2472 (
            .O(N__12447),
            .I(N__12442));
    LocalMux I__2471 (
            .O(N__12442),
            .I(N__12439));
    Span4Mux_h I__2470 (
            .O(N__12439),
            .I(N__12433));
    InMux I__2469 (
            .O(N__12438),
            .I(N__12430));
    InMux I__2468 (
            .O(N__12437),
            .I(N__12425));
    InMux I__2467 (
            .O(N__12436),
            .I(N__12425));
    Odrv4 I__2466 (
            .O(N__12433),
            .I(if_generate_plus_mult1_un68_sum_axbxc5));
    LocalMux I__2465 (
            .O(N__12430),
            .I(if_generate_plus_mult1_un68_sum_axbxc5));
    LocalMux I__2464 (
            .O(N__12425),
            .I(if_generate_plus_mult1_un68_sum_axbxc5));
    CascadeMux I__2463 (
            .O(N__12418),
            .I(N__12414));
    CascadeMux I__2462 (
            .O(N__12417),
            .I(N__12411));
    InMux I__2461 (
            .O(N__12414),
            .I(N__12407));
    InMux I__2460 (
            .O(N__12411),
            .I(N__12401));
    InMux I__2459 (
            .O(N__12410),
            .I(N__12401));
    LocalMux I__2458 (
            .O(N__12407),
            .I(N__12398));
    InMux I__2457 (
            .O(N__12406),
            .I(N__12395));
    LocalMux I__2456 (
            .O(N__12401),
            .I(N__12392));
    Span4Mux_h I__2455 (
            .O(N__12398),
            .I(N__12389));
    LocalMux I__2454 (
            .O(N__12395),
            .I(N__12386));
    Span4Mux_h I__2453 (
            .O(N__12392),
            .I(N__12383));
    Odrv4 I__2452 (
            .O(N__12389),
            .I(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2));
    Odrv4 I__2451 (
            .O(N__12386),
            .I(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2));
    Odrv4 I__2450 (
            .O(N__12383),
            .I(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2));
    InMux I__2449 (
            .O(N__12376),
            .I(N__12373));
    LocalMux I__2448 (
            .O(N__12373),
            .I(un114_pixel_1_0_3__un4_row_8Z0Z_7));
    InMux I__2447 (
            .O(N__12370),
            .I(N__12367));
    LocalMux I__2446 (
            .O(N__12367),
            .I(un114_pixel_1_0_3__un4_rowZ0Z_8));
    InMux I__2445 (
            .O(N__12364),
            .I(N__12361));
    LocalMux I__2444 (
            .O(N__12361),
            .I(N__12357));
    InMux I__2443 (
            .O(N__12360),
            .I(N__12354));
    Span4Mux_h I__2442 (
            .O(N__12357),
            .I(N__12351));
    LocalMux I__2441 (
            .O(N__12354),
            .I(N__12348));
    Odrv4 I__2440 (
            .O(N__12351),
            .I(row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1));
    Odrv12 I__2439 (
            .O(N__12348),
            .I(row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1));
    InMux I__2438 (
            .O(N__12343),
            .I(N__12339));
    InMux I__2437 (
            .O(N__12342),
            .I(N__12336));
    LocalMux I__2436 (
            .O(N__12339),
            .I(N__12333));
    LocalMux I__2435 (
            .O(N__12336),
            .I(N__12330));
    Span4Mux_v I__2434 (
            .O(N__12333),
            .I(N__12325));
    Span4Mux_h I__2433 (
            .O(N__12330),
            .I(N__12325));
    Odrv4 I__2432 (
            .O(N__12325),
            .I(row_1_if_generate_plus_mult1_un82_sum_c5));
    CascadeMux I__2431 (
            .O(N__12322),
            .I(un114_pixel_1_0_3__un4_rowZ0Z_8_cascade_));
    InMux I__2430 (
            .O(N__12319),
            .I(N__12316));
    LocalMux I__2429 (
            .O(N__12316),
            .I(N__12313));
    Odrv12 I__2428 (
            .O(N__12313),
            .I(un114_pixel_1_0_3__Pixel_3_sqmuxaZ0Z_0));
    InMux I__2427 (
            .O(N__12310),
            .I(N__12307));
    LocalMux I__2426 (
            .O(N__12307),
            .I(N__12303));
    InMux I__2425 (
            .O(N__12306),
            .I(N__12300));
    Odrv4 I__2424 (
            .O(N__12303),
            .I(Pixel_3_sqmuxa));
    LocalMux I__2423 (
            .O(N__12300),
            .I(Pixel_3_sqmuxa));
    InMux I__2422 (
            .O(N__12295),
            .I(charx_if_generate_plus_mult1_un75_sum_cry_1));
    InMux I__2421 (
            .O(N__12292),
            .I(N__12288));
    InMux I__2420 (
            .O(N__12291),
            .I(N__12285));
    LocalMux I__2419 (
            .O(N__12288),
            .I(N__12282));
    LocalMux I__2418 (
            .O(N__12285),
            .I(N__12275));
    Span4Mux_h I__2417 (
            .O(N__12282),
            .I(N__12275));
    InMux I__2416 (
            .O(N__12281),
            .I(N__12270));
    InMux I__2415 (
            .O(N__12280),
            .I(N__12270));
    Odrv4 I__2414 (
            .O(N__12275),
            .I(beamY_RNIHHB5F01Z0Z_4));
    LocalMux I__2413 (
            .O(N__12270),
            .I(beamY_RNIHHB5F01Z0Z_4));
    InMux I__2412 (
            .O(N__12265),
            .I(N__12260));
    InMux I__2411 (
            .O(N__12264),
            .I(N__12255));
    InMux I__2410 (
            .O(N__12263),
            .I(N__12255));
    LocalMux I__2409 (
            .O(N__12260),
            .I(N__12242));
    LocalMux I__2408 (
            .O(N__12255),
            .I(N__12239));
    InMux I__2407 (
            .O(N__12254),
            .I(N__12234));
    InMux I__2406 (
            .O(N__12253),
            .I(N__12234));
    InMux I__2405 (
            .O(N__12252),
            .I(N__12231));
    InMux I__2404 (
            .O(N__12251),
            .I(N__12228));
    InMux I__2403 (
            .O(N__12250),
            .I(N__12225));
    InMux I__2402 (
            .O(N__12249),
            .I(N__12222));
    InMux I__2401 (
            .O(N__12248),
            .I(N__12217));
    InMux I__2400 (
            .O(N__12247),
            .I(N__12217));
    InMux I__2399 (
            .O(N__12246),
            .I(N__12212));
    InMux I__2398 (
            .O(N__12245),
            .I(N__12209));
    Span4Mux_v I__2397 (
            .O(N__12242),
            .I(N__12203));
    Span4Mux_v I__2396 (
            .O(N__12239),
            .I(N__12203));
    LocalMux I__2395 (
            .O(N__12234),
            .I(N__12196));
    LocalMux I__2394 (
            .O(N__12231),
            .I(N__12196));
    LocalMux I__2393 (
            .O(N__12228),
            .I(N__12196));
    LocalMux I__2392 (
            .O(N__12225),
            .I(N__12189));
    LocalMux I__2391 (
            .O(N__12222),
            .I(N__12189));
    LocalMux I__2390 (
            .O(N__12217),
            .I(N__12189));
    InMux I__2389 (
            .O(N__12216),
            .I(N__12184));
    InMux I__2388 (
            .O(N__12215),
            .I(N__12184));
    LocalMux I__2387 (
            .O(N__12212),
            .I(N__12179));
    LocalMux I__2386 (
            .O(N__12209),
            .I(N__12179));
    InMux I__2385 (
            .O(N__12208),
            .I(N__12174));
    Span4Mux_h I__2384 (
            .O(N__12203),
            .I(N__12171));
    Span4Mux_v I__2383 (
            .O(N__12196),
            .I(N__12164));
    Span4Mux_v I__2382 (
            .O(N__12189),
            .I(N__12164));
    LocalMux I__2381 (
            .O(N__12184),
            .I(N__12164));
    Span4Mux_v I__2380 (
            .O(N__12179),
            .I(N__12161));
    InMux I__2379 (
            .O(N__12178),
            .I(N__12156));
    InMux I__2378 (
            .O(N__12177),
            .I(N__12156));
    LocalMux I__2377 (
            .O(N__12174),
            .I(beamYZ0Z_2));
    Odrv4 I__2376 (
            .O(N__12171),
            .I(beamYZ0Z_2));
    Odrv4 I__2375 (
            .O(N__12164),
            .I(beamYZ0Z_2));
    Odrv4 I__2374 (
            .O(N__12161),
            .I(beamYZ0Z_2));
    LocalMux I__2373 (
            .O(N__12156),
            .I(beamYZ0Z_2));
    CascadeMux I__2372 (
            .O(N__12145),
            .I(N__12142));
    InMux I__2371 (
            .O(N__12142),
            .I(N__12139));
    LocalMux I__2370 (
            .O(N__12139),
            .I(beamY_RNI7OE17CZ0Z_0));
    InMux I__2369 (
            .O(N__12136),
            .I(N__12133));
    LocalMux I__2368 (
            .O(N__12133),
            .I(N__12130));
    Odrv4 I__2367 (
            .O(N__12130),
            .I(beamY_RNIVU1O9RZ0Z_1));
    InMux I__2366 (
            .O(N__12127),
            .I(N__12124));
    LocalMux I__2365 (
            .O(N__12124),
            .I(font_un126_pixel_6_bm));
    CascadeMux I__2364 (
            .O(N__12121),
            .I(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_));
    InMux I__2363 (
            .O(N__12118),
            .I(N__12114));
    InMux I__2362 (
            .O(N__12117),
            .I(N__12111));
    LocalMux I__2361 (
            .O(N__12114),
            .I(N__12108));
    LocalMux I__2360 (
            .O(N__12111),
            .I(N__12105));
    Span4Mux_v I__2359 (
            .O(N__12108),
            .I(N__12102));
    Span4Mux_h I__2358 (
            .O(N__12105),
            .I(N__12099));
    Odrv4 I__2357 (
            .O(N__12102),
            .I(un15_beamy));
    Odrv4 I__2356 (
            .O(N__12099),
            .I(un15_beamy));
    CascadeMux I__2355 (
            .O(N__12094),
            .I(r_i1_mux_cascade_));
    CascadeMux I__2354 (
            .O(N__12091),
            .I(un114_pixel_1_0_3__font_un126_pixel_mZ0Z_1_cascade_));
    InMux I__2353 (
            .O(N__12088),
            .I(N__12085));
    LocalMux I__2352 (
            .O(N__12085),
            .I(N__12082));
    Span4Mux_v I__2351 (
            .O(N__12082),
            .I(N__12079));
    Odrv4 I__2350 (
            .O(N__12079),
            .I(chary_24));
    CascadeMux I__2349 (
            .O(N__12076),
            .I(un114_pixel_1_0_3__font_un126_pixel_m_1_0_cascade_));
    InMux I__2348 (
            .O(N__12073),
            .I(N__12070));
    LocalMux I__2347 (
            .O(N__12070),
            .I(chary_23));
    InMux I__2346 (
            .O(N__12067),
            .I(N__12064));
    LocalMux I__2345 (
            .O(N__12064),
            .I(un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3));
    InMux I__2344 (
            .O(N__12061),
            .I(N__12057));
    InMux I__2343 (
            .O(N__12060),
            .I(N__12054));
    LocalMux I__2342 (
            .O(N__12057),
            .I(N__12051));
    LocalMux I__2341 (
            .O(N__12054),
            .I(N__12048));
    Span4Mux_h I__2340 (
            .O(N__12051),
            .I(N__12045));
    Span12Mux_s5_v I__2339 (
            .O(N__12048),
            .I(N__12042));
    Span4Mux_h I__2338 (
            .O(N__12045),
            .I(N__12039));
    Odrv12 I__2337 (
            .O(N__12042),
            .I(un1_beamylto9));
    Odrv4 I__2336 (
            .O(N__12039),
            .I(un1_beamylto9));
    CascadeMux I__2335 (
            .O(N__12034),
            .I(un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3_cascade_));
    InMux I__2334 (
            .O(N__12031),
            .I(N__12028));
    LocalMux I__2333 (
            .O(N__12028),
            .I(Pixel_r_sn));
    CascadeMux I__2332 (
            .O(N__12025),
            .I(N__12020));
    CascadeMux I__2331 (
            .O(N__12024),
            .I(N__12015));
    InMux I__2330 (
            .O(N__12023),
            .I(N__12012));
    InMux I__2329 (
            .O(N__12020),
            .I(N__12009));
    InMux I__2328 (
            .O(N__12019),
            .I(N__12004));
    InMux I__2327 (
            .O(N__12018),
            .I(N__12004));
    InMux I__2326 (
            .O(N__12015),
            .I(N__11999));
    LocalMux I__2325 (
            .O(N__12012),
            .I(N__11994));
    LocalMux I__2324 (
            .O(N__12009),
            .I(N__11994));
    LocalMux I__2323 (
            .O(N__12004),
            .I(N__11991));
    CascadeMux I__2322 (
            .O(N__12003),
            .I(N__11985));
    InMux I__2321 (
            .O(N__12002),
            .I(N__11982));
    LocalMux I__2320 (
            .O(N__11999),
            .I(N__11979));
    Span4Mux_h I__2319 (
            .O(N__11994),
            .I(N__11976));
    Span4Mux_h I__2318 (
            .O(N__11991),
            .I(N__11973));
    InMux I__2317 (
            .O(N__11990),
            .I(N__11966));
    InMux I__2316 (
            .O(N__11989),
            .I(N__11966));
    InMux I__2315 (
            .O(N__11988),
            .I(N__11966));
    InMux I__2314 (
            .O(N__11985),
            .I(N__11963));
    LocalMux I__2313 (
            .O(N__11982),
            .I(beamXZ0Z_0));
    Odrv4 I__2312 (
            .O(N__11979),
            .I(beamXZ0Z_0));
    Odrv4 I__2311 (
            .O(N__11976),
            .I(beamXZ0Z_0));
    Odrv4 I__2310 (
            .O(N__11973),
            .I(beamXZ0Z_0));
    LocalMux I__2309 (
            .O(N__11966),
            .I(beamXZ0Z_0));
    LocalMux I__2308 (
            .O(N__11963),
            .I(beamXZ0Z_0));
    CascadeMux I__2307 (
            .O(N__11950),
            .I(N_364_cascade_));
    CascadeMux I__2306 (
            .O(N__11947),
            .I(un116_pixel_7_ns_1_4_cascade_));
    InMux I__2305 (
            .O(N__11944),
            .I(N__11941));
    LocalMux I__2304 (
            .O(N__11941),
            .I(beamY_RNI2L0T663Z0Z_0));
    InMux I__2303 (
            .O(N__11938),
            .I(N__11935));
    LocalMux I__2302 (
            .O(N__11935),
            .I(column_0111_1_0));
    InMux I__2301 (
            .O(N__11932),
            .I(N__11929));
    LocalMux I__2300 (
            .O(N__11929),
            .I(beamY_RNI1J75181Z0Z_1));
    CascadeMux I__2299 (
            .O(N__11926),
            .I(font_un126_pixel_6_am_cascade_));
    InMux I__2298 (
            .O(N__11923),
            .I(N__11920));
    LocalMux I__2297 (
            .O(N__11920),
            .I(N__11917));
    Span4Mux_h I__2296 (
            .O(N__11917),
            .I(N__11914));
    Odrv4 I__2295 (
            .O(N__11914),
            .I(un1_beamy_0));
    CascadeMux I__2294 (
            .O(N__11911),
            .I(N_1075_0_cascade_));
    InMux I__2293 (
            .O(N__11908),
            .I(N__11905));
    LocalMux I__2292 (
            .O(N__11905),
            .I(N__11902));
    Odrv4 I__2291 (
            .O(N__11902),
            .I(N_400));
    CascadeMux I__2290 (
            .O(N__11899),
            .I(Pixel_r_rn_0_cascade_));
    IoInMux I__2289 (
            .O(N__11896),
            .I(N__11893));
    LocalMux I__2288 (
            .O(N__11893),
            .I(N__11890));
    Span4Mux_s3_v I__2287 (
            .O(N__11890),
            .I(N__11887));
    Odrv4 I__2286 (
            .O(N__11887),
            .I(Pixel_c));
    ClkMux I__2285 (
            .O(N__11884),
            .I(N__11845));
    ClkMux I__2284 (
            .O(N__11883),
            .I(N__11845));
    ClkMux I__2283 (
            .O(N__11882),
            .I(N__11845));
    ClkMux I__2282 (
            .O(N__11881),
            .I(N__11845));
    ClkMux I__2281 (
            .O(N__11880),
            .I(N__11845));
    ClkMux I__2280 (
            .O(N__11879),
            .I(N__11845));
    ClkMux I__2279 (
            .O(N__11878),
            .I(N__11845));
    ClkMux I__2278 (
            .O(N__11877),
            .I(N__11845));
    ClkMux I__2277 (
            .O(N__11876),
            .I(N__11845));
    ClkMux I__2276 (
            .O(N__11875),
            .I(N__11845));
    ClkMux I__2275 (
            .O(N__11874),
            .I(N__11845));
    ClkMux I__2274 (
            .O(N__11873),
            .I(N__11845));
    ClkMux I__2273 (
            .O(N__11872),
            .I(N__11845));
    GlobalMux I__2272 (
            .O(N__11845),
            .I(N__11842));
    gio2CtrlBuf I__2271 (
            .O(N__11842),
            .I(PixelClock_g));
    InMux I__2270 (
            .O(N__11839),
            .I(N__11836));
    LocalMux I__2269 (
            .O(N__11836),
            .I(N__11833));
    Span4Mux_v I__2268 (
            .O(N__11833),
            .I(N__11830));
    Odrv4 I__2267 (
            .O(N__11830),
            .I(font_un28_pixel_0_0_29));
    InMux I__2266 (
            .O(N__11827),
            .I(N__11824));
    LocalMux I__2265 (
            .O(N__11824),
            .I(font_un126_pixel_2_bm));
    InMux I__2264 (
            .O(N__11821),
            .I(N__11818));
    LocalMux I__2263 (
            .O(N__11818),
            .I(un114_pixel_1_0_3__font_un126_pixel_7_d_ns_1_0_0));
    CascadeMux I__2262 (
            .O(N__11815),
            .I(font_un3_pixel_29_cascade_));
    InMux I__2261 (
            .O(N__11812),
            .I(N__11809));
    LocalMux I__2260 (
            .O(N__11809),
            .I(un116_pixel_5_bm_6));
    InMux I__2259 (
            .O(N__11806),
            .I(N__11803));
    LocalMux I__2258 (
            .O(N__11803),
            .I(un116_pixel_4_bm_1));
    CascadeMux I__2257 (
            .O(N__11800),
            .I(beamY_RNI1C50FS3Z0Z_0_cascade_));
    CascadeMux I__2256 (
            .O(N__11797),
            .I(un116_pixel_3_bm_1_6_cascade_));
    InMux I__2255 (
            .O(N__11794),
            .I(N__11788));
    InMux I__2254 (
            .O(N__11793),
            .I(N__11788));
    LocalMux I__2253 (
            .O(N__11788),
            .I(N__11785));
    Odrv4 I__2252 (
            .O(N__11785),
            .I(beamY_RNIOHI2NGZ0Z_0));
    CascadeMux I__2251 (
            .O(N__11782),
            .I(N_1556_0_cascade_));
    InMux I__2250 (
            .O(N__11779),
            .I(N__11776));
    LocalMux I__2249 (
            .O(N__11776),
            .I(N__11773));
    Odrv4 I__2248 (
            .O(N__11773),
            .I(N_347_0));
    CascadeMux I__2247 (
            .O(N__11770),
            .I(N__11767));
    InMux I__2246 (
            .O(N__11767),
            .I(N__11764));
    LocalMux I__2245 (
            .O(N__11764),
            .I(font_un28_pixel_0_29));
    InMux I__2244 (
            .O(N__11761),
            .I(N__11758));
    LocalMux I__2243 (
            .O(N__11758),
            .I(N_368_0));
    CascadeMux I__2242 (
            .O(N__11755),
            .I(un114_pixel_1_0_3__font_un126_pixel_1_d_ns_1_0_cascade_));
    InMux I__2241 (
            .O(N__11752),
            .I(N__11749));
    LocalMux I__2240 (
            .O(N__11749),
            .I(N_389_0));
    InMux I__2239 (
            .O(N__11746),
            .I(N__11743));
    LocalMux I__2238 (
            .O(N__11743),
            .I(N_346_0_0_1));
    CascadeMux I__2237 (
            .O(N__11740),
            .I(g0_cascade_));
    CascadeMux I__2236 (
            .O(N__11737),
            .I(N_36_cascade_));
    CascadeMux I__2235 (
            .O(N__11734),
            .I(un116_pixel_3_ns_1_1_cascade_));
    InMux I__2234 (
            .O(N__11731),
            .I(N__11728));
    LocalMux I__2233 (
            .O(N__11728),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLMZ0Z67));
    InMux I__2232 (
            .O(N__11725),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__2231 (
            .O(N__11722),
            .I(N__11719));
    LocalMux I__2230 (
            .O(N__11719),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSAZ0));
    InMux I__2229 (
            .O(N__11716),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__2228 (
            .O(N__11713),
            .I(N__11710));
    LocalMux I__2227 (
            .O(N__11710),
            .I(charx_if_generate_plus_mult1_un61_sum_axb_5));
    InMux I__2226 (
            .O(N__11707),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__2225 (
            .O(N__11704),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0_cascade_));
    CascadeMux I__2224 (
            .O(N__11701),
            .I(N__11697));
    InMux I__2223 (
            .O(N__11700),
            .I(N__11693));
    InMux I__2222 (
            .O(N__11697),
            .I(N__11688));
    InMux I__2221 (
            .O(N__11696),
            .I(N__11688));
    LocalMux I__2220 (
            .O(N__11693),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0));
    LocalMux I__2219 (
            .O(N__11688),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0));
    CascadeMux I__2218 (
            .O(N__11683),
            .I(N__11679));
    CascadeMux I__2217 (
            .O(N__11682),
            .I(N__11676));
    InMux I__2216 (
            .O(N__11679),
            .I(N__11671));
    InMux I__2215 (
            .O(N__11676),
            .I(N__11671));
    LocalMux I__2214 (
            .O(N__11671),
            .I(charx_if_generate_plus_mult1_un54_sum_i_5));
    IoInMux I__2213 (
            .O(N__11668),
            .I(N__11665));
    LocalMux I__2212 (
            .O(N__11665),
            .I(VSync_c));
    InMux I__2211 (
            .O(N__11662),
            .I(N__11659));
    LocalMux I__2210 (
            .O(N__11659),
            .I(un116_pixel_3_am_2));
    InMux I__2209 (
            .O(N__11656),
            .I(N__11653));
    LocalMux I__2208 (
            .O(N__11653),
            .I(N__11646));
    InMux I__2207 (
            .O(N__11652),
            .I(N__11642));
    InMux I__2206 (
            .O(N__11651),
            .I(N__11637));
    InMux I__2205 (
            .O(N__11650),
            .I(N__11637));
    InMux I__2204 (
            .O(N__11649),
            .I(N__11634));
    Span4Mux_v I__2203 (
            .O(N__11646),
            .I(N__11631));
    InMux I__2202 (
            .O(N__11645),
            .I(N__11628));
    LocalMux I__2201 (
            .O(N__11642),
            .I(N__11623));
    LocalMux I__2200 (
            .O(N__11637),
            .I(N__11623));
    LocalMux I__2199 (
            .O(N__11634),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__2198 (
            .O(N__11631),
            .I(charx_if_generate_plus_mult1_un47_sum));
    LocalMux I__2197 (
            .O(N__11628),
            .I(charx_if_generate_plus_mult1_un47_sum));
    Odrv4 I__2196 (
            .O(N__11623),
            .I(charx_if_generate_plus_mult1_un47_sum));
    InMux I__2195 (
            .O(N__11614),
            .I(N__11611));
    LocalMux I__2194 (
            .O(N__11611),
            .I(charx_if_generate_plus_mult1_un47_sum_i));
    InMux I__2193 (
            .O(N__11608),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__2192 (
            .O(N__11605),
            .I(N__11601));
    InMux I__2191 (
            .O(N__11604),
            .I(N__11598));
    LocalMux I__2190 (
            .O(N__11601),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6));
    LocalMux I__2189 (
            .O(N__11598),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6));
    CascadeMux I__2188 (
            .O(N__11593),
            .I(N__11590));
    InMux I__2187 (
            .O(N__11590),
            .I(N__11587));
    LocalMux I__2186 (
            .O(N__11587),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0OZ0Z3));
    InMux I__2185 (
            .O(N__11584),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__2184 (
            .O(N__11581),
            .I(N__11578));
    LocalMux I__2183 (
            .O(N__11578),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCDZ0Z16));
    CascadeMux I__2182 (
            .O(N__11575),
            .I(N__11571));
    CascadeMux I__2181 (
            .O(N__11574),
            .I(N__11568));
    InMux I__2180 (
            .O(N__11571),
            .I(N__11563));
    InMux I__2179 (
            .O(N__11568),
            .I(N__11563));
    LocalMux I__2178 (
            .O(N__11563),
            .I(charx_if_generate_plus_mult1_un47_sum_i_5));
    InMux I__2177 (
            .O(N__11560),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__2176 (
            .O(N__11557),
            .I(N__11554));
    LocalMux I__2175 (
            .O(N__11554),
            .I(charx_if_generate_plus_mult1_un54_sum_axb_5));
    InMux I__2174 (
            .O(N__11551),
            .I(charx_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__2173 (
            .O(N__11548),
            .I(N__11539));
    InMux I__2172 (
            .O(N__11547),
            .I(N__11539));
    InMux I__2171 (
            .O(N__11546),
            .I(N__11532));
    InMux I__2170 (
            .O(N__11545),
            .I(N__11532));
    InMux I__2169 (
            .O(N__11544),
            .I(N__11529));
    LocalMux I__2168 (
            .O(N__11539),
            .I(N__11526));
    InMux I__2167 (
            .O(N__11538),
            .I(N__11523));
    InMux I__2166 (
            .O(N__11537),
            .I(N__11520));
    LocalMux I__2165 (
            .O(N__11532),
            .I(N__11517));
    LocalMux I__2164 (
            .O(N__11529),
            .I(N__11514));
    Span4Mux_v I__2163 (
            .O(N__11526),
            .I(N__11511));
    LocalMux I__2162 (
            .O(N__11523),
            .I(N__11506));
    LocalMux I__2161 (
            .O(N__11520),
            .I(N__11506));
    Span4Mux_s3_v I__2160 (
            .O(N__11517),
            .I(N__11503));
    Odrv12 I__2159 (
            .O(N__11514),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv4 I__2158 (
            .O(N__11511),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv4 I__2157 (
            .O(N__11506),
            .I(charx_if_generate_plus_mult1_un54_sum));
    Odrv4 I__2156 (
            .O(N__11503),
            .I(charx_if_generate_plus_mult1_un54_sum));
    InMux I__2155 (
            .O(N__11494),
            .I(N__11491));
    LocalMux I__2154 (
            .O(N__11491),
            .I(charx_if_generate_plus_mult1_un54_sum_i));
    InMux I__2153 (
            .O(N__11488),
            .I(charx_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__2152 (
            .O(N__11485),
            .I(N__11482));
    LocalMux I__2151 (
            .O(N__11482),
            .I(column_1_if_generate_plus_mult1_un47_sum0_3));
    CascadeMux I__2150 (
            .O(N__11479),
            .I(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_));
    InMux I__2149 (
            .O(N__11476),
            .I(N__11473));
    LocalMux I__2148 (
            .O(N__11473),
            .I(if_generate_plus_mult1_un54_sum_axb_4_l_fx));
    InMux I__2147 (
            .O(N__11470),
            .I(N__11467));
    LocalMux I__2146 (
            .O(N__11467),
            .I(N__11464));
    Odrv4 I__2145 (
            .O(N__11464),
            .I(charx_if_generate_plus_mult1_un40_sum_i));
    InMux I__2144 (
            .O(N__11461),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_1));
    InMux I__2143 (
            .O(N__11458),
            .I(N__11453));
    InMux I__2142 (
            .O(N__11457),
            .I(N__11450));
    InMux I__2141 (
            .O(N__11456),
            .I(N__11447));
    LocalMux I__2140 (
            .O(N__11453),
            .I(N__11442));
    LocalMux I__2139 (
            .O(N__11450),
            .I(N__11442));
    LocalMux I__2138 (
            .O(N__11447),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3));
    Odrv4 I__2137 (
            .O(N__11442),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3));
    CascadeMux I__2136 (
            .O(N__11437),
            .I(N__11434));
    InMux I__2135 (
            .O(N__11434),
            .I(N__11431));
    LocalMux I__2134 (
            .O(N__11431),
            .I(N__11428));
    Odrv12 I__2133 (
            .O(N__11428),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEBZ0Z2));
    InMux I__2132 (
            .O(N__11425),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__2131 (
            .O(N__11422),
            .I(N__11419));
    LocalMux I__2130 (
            .O(N__11419),
            .I(N__11416));
    Odrv4 I__2129 (
            .O(N__11416),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLITZ0Z2));
    CascadeMux I__2128 (
            .O(N__11413),
            .I(N__11409));
    CascadeMux I__2127 (
            .O(N__11412),
            .I(N__11406));
    InMux I__2126 (
            .O(N__11409),
            .I(N__11401));
    InMux I__2125 (
            .O(N__11406),
            .I(N__11401));
    LocalMux I__2124 (
            .O(N__11401),
            .I(charx_if_generate_plus_mult1_un40_sum_i_5));
    InMux I__2123 (
            .O(N__11398),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__2122 (
            .O(N__11395),
            .I(N__11392));
    LocalMux I__2121 (
            .O(N__11392),
            .I(N__11389));
    Odrv4 I__2120 (
            .O(N__11389),
            .I(charx_if_generate_plus_mult1_un47_sum_axb_5));
    InMux I__2119 (
            .O(N__11386),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__2118 (
            .O(N__11383),
            .I(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6_cascade_));
    CascadeMux I__2117 (
            .O(N__11380),
            .I(N__11377));
    InMux I__2116 (
            .O(N__11377),
            .I(N__11374));
    LocalMux I__2115 (
            .O(N__11374),
            .I(un5_visiblex_i_25));
    CascadeMux I__2114 (
            .O(N__11371),
            .I(N__11368));
    InMux I__2113 (
            .O(N__11368),
            .I(N__11365));
    LocalMux I__2112 (
            .O(N__11365),
            .I(if_generate_plus_mult1_un47_sum_0_cry_3_ma));
    CascadeMux I__2111 (
            .O(N__11362),
            .I(N__11359));
    InMux I__2110 (
            .O(N__11359),
            .I(N__11356));
    LocalMux I__2109 (
            .O(N__11356),
            .I(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx));
    InMux I__2108 (
            .O(N__11353),
            .I(N__11350));
    LocalMux I__2107 (
            .O(N__11350),
            .I(N__11347));
    Span4Mux_h I__2106 (
            .O(N__11347),
            .I(N__11344));
    Odrv4 I__2105 (
            .O(N__11344),
            .I(if_generate_plus_mult1_un54_sum_cry_2_s));
    InMux I__2104 (
            .O(N__11341),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_1));
    CascadeMux I__2103 (
            .O(N__11338),
            .I(N__11335));
    InMux I__2102 (
            .O(N__11335),
            .I(N__11332));
    LocalMux I__2101 (
            .O(N__11332),
            .I(N__11329));
    Span4Mux_h I__2100 (
            .O(N__11329),
            .I(N__11326));
    Odrv4 I__2099 (
            .O(N__11326),
            .I(if_generate_plus_mult1_un54_sum_cry_3_s));
    InMux I__2098 (
            .O(N__11323),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__2097 (
            .O(N__11320),
            .I(N__11317));
    LocalMux I__2096 (
            .O(N__11317),
            .I(N__11314));
    Odrv12 I__2095 (
            .O(N__11314),
            .I(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5));
    InMux I__2094 (
            .O(N__11311),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__2093 (
            .O(N__11308),
            .I(column_1_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__2092 (
            .O(N__11305),
            .I(N__11302));
    LocalMux I__2091 (
            .O(N__11302),
            .I(charx_if_generate_plus_mult1_un40_sum_axb_5));
    InMux I__2090 (
            .O(N__11299),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__2089 (
            .O(N__11296),
            .I(N__11293));
    LocalMux I__2088 (
            .O(N__11293),
            .I(charx_if_generate_plus_mult1_un33_sum_i));
    InMux I__2087 (
            .O(N__11290),
            .I(N__11287));
    LocalMux I__2086 (
            .O(N__11287),
            .I(charx_if_generate_plus_mult1_un26_sum_i));
    InMux I__2085 (
            .O(N__11284),
            .I(N__11281));
    LocalMux I__2084 (
            .O(N__11281),
            .I(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx));
    InMux I__2083 (
            .O(N__11278),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_1));
    InMux I__2082 (
            .O(N__11275),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_2));
    InMux I__2081 (
            .O(N__11272),
            .I(N__11269));
    LocalMux I__2080 (
            .O(N__11269),
            .I(N__11266));
    Odrv4 I__2079 (
            .O(N__11266),
            .I(N_204_0_i));
    InMux I__2078 (
            .O(N__11263),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_3));
    InMux I__2077 (
            .O(N__11260),
            .I(column_1_if_generate_plus_mult1_un47_sum_0_cry_4));
    InMux I__2076 (
            .O(N__11257),
            .I(N__11254));
    LocalMux I__2075 (
            .O(N__11254),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328));
    InMux I__2074 (
            .O(N__11251),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__2073 (
            .O(N__11248),
            .I(N__11245));
    LocalMux I__2072 (
            .O(N__11245),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HLZ0));
    InMux I__2071 (
            .O(N__11242),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__2070 (
            .O(N__11239),
            .I(N__11236));
    LocalMux I__2069 (
            .O(N__11236),
            .I(charx_if_generate_plus_mult1_un33_sum_axb_5));
    InMux I__2068 (
            .O(N__11233),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4));
    CascadeMux I__2067 (
            .O(N__11230),
            .I(N__11226));
    InMux I__2066 (
            .O(N__11229),
            .I(N__11222));
    InMux I__2065 (
            .O(N__11226),
            .I(N__11217));
    InMux I__2064 (
            .O(N__11225),
            .I(N__11217));
    LocalMux I__2063 (
            .O(N__11222),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5));
    LocalMux I__2062 (
            .O(N__11217),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5));
    CascadeMux I__2061 (
            .O(N__11212),
            .I(N__11208));
    CascadeMux I__2060 (
            .O(N__11211),
            .I(N__11205));
    InMux I__2059 (
            .O(N__11208),
            .I(N__11200));
    InMux I__2058 (
            .O(N__11205),
            .I(N__11200));
    LocalMux I__2057 (
            .O(N__11200),
            .I(charx_if_generate_plus_mult1_un26_sum_i_5));
    InMux I__2056 (
            .O(N__11197),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_1));
    InMux I__2055 (
            .O(N__11194),
            .I(N__11189));
    InMux I__2054 (
            .O(N__11193),
            .I(N__11186));
    InMux I__2053 (
            .O(N__11192),
            .I(N__11183));
    LocalMux I__2052 (
            .O(N__11189),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072));
    LocalMux I__2051 (
            .O(N__11186),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072));
    LocalMux I__2050 (
            .O(N__11183),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072));
    CascadeMux I__2049 (
            .O(N__11176),
            .I(N__11173));
    InMux I__2048 (
            .O(N__11173),
            .I(N__11170));
    LocalMux I__2047 (
            .O(N__11170),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0));
    InMux I__2046 (
            .O(N__11167),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__2045 (
            .O(N__11164),
            .I(N__11161));
    LocalMux I__2044 (
            .O(N__11161),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0));
    CascadeMux I__2043 (
            .O(N__11158),
            .I(N__11154));
    CascadeMux I__2042 (
            .O(N__11157),
            .I(N__11151));
    InMux I__2041 (
            .O(N__11154),
            .I(N__11146));
    InMux I__2040 (
            .O(N__11151),
            .I(N__11146));
    LocalMux I__2039 (
            .O(N__11146),
            .I(charx_if_generate_plus_mult1_un33_sum_i_5));
    InMux I__2038 (
            .O(N__11143),
            .I(charx_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__2037 (
            .O(N__11140),
            .I(N__11134));
    InMux I__2036 (
            .O(N__11139),
            .I(N__11134));
    LocalMux I__2035 (
            .O(N__11134),
            .I(un5_rowlto3_i));
    InMux I__2034 (
            .O(N__11131),
            .I(N__11128));
    LocalMux I__2033 (
            .O(N__11128),
            .I(N_575_i));
    InMux I__2032 (
            .O(N__11125),
            .I(N__11122));
    LocalMux I__2031 (
            .O(N__11122),
            .I(if_generate_plus_mult1_un61_sum_cry_2_s));
    InMux I__2030 (
            .O(N__11119),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_1));
    CascadeMux I__2029 (
            .O(N__11116),
            .I(N__11113));
    InMux I__2028 (
            .O(N__11113),
            .I(N__11110));
    LocalMux I__2027 (
            .O(N__11110),
            .I(if_generate_plus_mult1_un61_sum_cry_3_s));
    InMux I__2026 (
            .O(N__11107),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__2025 (
            .O(N__11104),
            .I(N__11101));
    LocalMux I__2024 (
            .O(N__11101),
            .I(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5));
    InMux I__2023 (
            .O(N__11098),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__2022 (
            .O(N__11095),
            .I(column_1_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__2021 (
            .O(N__11092),
            .I(N__11088));
    InMux I__2020 (
            .O(N__11091),
            .I(N__11085));
    InMux I__2019 (
            .O(N__11088),
            .I(N__11082));
    LocalMux I__2018 (
            .O(N__11085),
            .I(column_1_if_generate_plus_mult1_un54_sum_i_5));
    LocalMux I__2017 (
            .O(N__11082),
            .I(column_1_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__2016 (
            .O(N__11077),
            .I(charx_if_generate_plus_mult1_un33_sum_cry_1));
    InMux I__2015 (
            .O(N__11074),
            .I(N__11071));
    LocalMux I__2014 (
            .O(N__11071),
            .I(N_41));
    CEMux I__2013 (
            .O(N__11068),
            .I(N__11062));
    CEMux I__2012 (
            .O(N__11067),
            .I(N__11059));
    CEMux I__2011 (
            .O(N__11066),
            .I(N__11054));
    CEMux I__2010 (
            .O(N__11065),
            .I(N__11051));
    LocalMux I__2009 (
            .O(N__11062),
            .I(N__11046));
    LocalMux I__2008 (
            .O(N__11059),
            .I(N__11046));
    CEMux I__2007 (
            .O(N__11058),
            .I(N__11043));
    CEMux I__2006 (
            .O(N__11057),
            .I(N__11037));
    LocalMux I__2005 (
            .O(N__11054),
            .I(N__11032));
    LocalMux I__2004 (
            .O(N__11051),
            .I(N__11032));
    Span4Mux_v I__2003 (
            .O(N__11046),
            .I(N__11027));
    LocalMux I__2002 (
            .O(N__11043),
            .I(N__11027));
    InMux I__2001 (
            .O(N__11042),
            .I(N__11023));
    InMux I__2000 (
            .O(N__11041),
            .I(N__11020));
    InMux I__1999 (
            .O(N__11040),
            .I(N__11017));
    LocalMux I__1998 (
            .O(N__11037),
            .I(N__11010));
    Span4Mux_v I__1997 (
            .O(N__11032),
            .I(N__11010));
    Span4Mux_s1_h I__1996 (
            .O(N__11027),
            .I(N__11010));
    InMux I__1995 (
            .O(N__11026),
            .I(N__11007));
    LocalMux I__1994 (
            .O(N__11023),
            .I(N__11004));
    LocalMux I__1993 (
            .O(N__11020),
            .I(N__10999));
    LocalMux I__1992 (
            .O(N__11017),
            .I(N__10999));
    Span4Mux_h I__1991 (
            .O(N__11010),
            .I(N__10996));
    LocalMux I__1990 (
            .O(N__11007),
            .I(N__10993));
    Span4Mux_h I__1989 (
            .O(N__11004),
            .I(N__10990));
    Span4Mux_v I__1988 (
            .O(N__10999),
            .I(N__10985));
    Span4Mux_h I__1987 (
            .O(N__10996),
            .I(N__10985));
    Odrv4 I__1986 (
            .O(N__10993),
            .I(un3_beamx_0));
    Odrv4 I__1985 (
            .O(N__10990),
            .I(un3_beamx_0));
    Odrv4 I__1984 (
            .O(N__10985),
            .I(un3_beamx_0));
    InMux I__1983 (
            .O(N__10978),
            .I(N__10971));
    InMux I__1982 (
            .O(N__10977),
            .I(N__10967));
    InMux I__1981 (
            .O(N__10976),
            .I(N__10964));
    InMux I__1980 (
            .O(N__10975),
            .I(N__10959));
    InMux I__1979 (
            .O(N__10974),
            .I(N__10959));
    LocalMux I__1978 (
            .O(N__10971),
            .I(N__10956));
    InMux I__1977 (
            .O(N__10970),
            .I(N__10951));
    LocalMux I__1976 (
            .O(N__10967),
            .I(N__10948));
    LocalMux I__1975 (
            .O(N__10964),
            .I(N__10945));
    LocalMux I__1974 (
            .O(N__10959),
            .I(N__10942));
    Span4Mux_v I__1973 (
            .O(N__10956),
            .I(N__10939));
    InMux I__1972 (
            .O(N__10955),
            .I(N__10934));
    InMux I__1971 (
            .O(N__10954),
            .I(N__10934));
    LocalMux I__1970 (
            .O(N__10951),
            .I(N__10927));
    Span4Mux_v I__1969 (
            .O(N__10948),
            .I(N__10927));
    Span4Mux_v I__1968 (
            .O(N__10945),
            .I(N__10927));
    Span4Mux_s3_h I__1967 (
            .O(N__10942),
            .I(N__10924));
    Sp12to4 I__1966 (
            .O(N__10939),
            .I(N__10919));
    LocalMux I__1965 (
            .O(N__10934),
            .I(N__10919));
    Odrv4 I__1964 (
            .O(N__10927),
            .I(un5_beamx_0));
    Odrv4 I__1963 (
            .O(N__10924),
            .I(un5_beamx_0));
    Odrv12 I__1962 (
            .O(N__10919),
            .I(un5_beamx_0));
    InMux I__1961 (
            .O(N__10912),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_1));
    InMux I__1960 (
            .O(N__10909),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__1959 (
            .O(N__10906),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__1958 (
            .O(N__10903),
            .I(column_1_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1957 (
            .O(N__10900),
            .I(N__10897));
    InMux I__1956 (
            .O(N__10897),
            .I(N__10894));
    LocalMux I__1955 (
            .O(N__10894),
            .I(column_1_if_generate_plus_mult1_un61_sum_iZ0));
    InMux I__1954 (
            .O(N__10891),
            .I(N__10887));
    InMux I__1953 (
            .O(N__10890),
            .I(N__10884));
    LocalMux I__1952 (
            .O(N__10887),
            .I(N__10874));
    LocalMux I__1951 (
            .O(N__10884),
            .I(N__10871));
    InMux I__1950 (
            .O(N__10883),
            .I(N__10860));
    InMux I__1949 (
            .O(N__10882),
            .I(N__10860));
    InMux I__1948 (
            .O(N__10881),
            .I(N__10860));
    InMux I__1947 (
            .O(N__10880),
            .I(N__10860));
    InMux I__1946 (
            .O(N__10879),
            .I(N__10860));
    InMux I__1945 (
            .O(N__10878),
            .I(N__10855));
    InMux I__1944 (
            .O(N__10877),
            .I(N__10855));
    Span4Mux_s3_h I__1943 (
            .O(N__10874),
            .I(N__10852));
    Span4Mux_h I__1942 (
            .O(N__10871),
            .I(N__10847));
    LocalMux I__1941 (
            .O(N__10860),
            .I(N__10847));
    LocalMux I__1940 (
            .O(N__10855),
            .I(row_1_if_generate_plus_mult1_un54_sum_cZ0Z5));
    Odrv4 I__1939 (
            .O(N__10852),
            .I(row_1_if_generate_plus_mult1_un54_sum_cZ0Z5));
    Odrv4 I__1938 (
            .O(N__10847),
            .I(row_1_if_generate_plus_mult1_un54_sum_cZ0Z5));
    CascadeMux I__1937 (
            .O(N__10840),
            .I(un116_pixel_5_ns_1Z0Z_4_cascade_));
    InMux I__1936 (
            .O(N__10837),
            .I(N__10834));
    LocalMux I__1935 (
            .O(N__10834),
            .I(un116_pixel_5_ns_2));
    InMux I__1934 (
            .O(N__10831),
            .I(N__10828));
    LocalMux I__1933 (
            .O(N__10828),
            .I(N_362));
    CascadeMux I__1932 (
            .O(N__10825),
            .I(un116_pixel_7_ns_1_6_cascade_));
    InMux I__1931 (
            .O(N__10822),
            .I(N__10819));
    LocalMux I__1930 (
            .O(N__10819),
            .I(N_379));
    InMux I__1929 (
            .O(N__10816),
            .I(N__10813));
    LocalMux I__1928 (
            .O(N__10813),
            .I(N__10810));
    Odrv12 I__1927 (
            .O(N__10810),
            .I(un116_pixel_3_ns_2));
    CascadeMux I__1926 (
            .O(N__10807),
            .I(beamY_RNI57H3N31_0Z0Z_1_cascade_));
    InMux I__1925 (
            .O(N__10804),
            .I(N__10801));
    LocalMux I__1924 (
            .O(N__10801),
            .I(beamY_RNI896FQ3Z0Z_0));
    CascadeMux I__1923 (
            .O(N__10798),
            .I(beamY_RNI896FQ3Z0Z_0_cascade_));
    InMux I__1922 (
            .O(N__10795),
            .I(N__10792));
    LocalMux I__1921 (
            .O(N__10792),
            .I(beamY_RNI57H3N31Z0Z_1));
    CascadeMux I__1920 (
            .O(N__10789),
            .I(un116_pixel_2_ns_1_0_6_cascade_));
    InMux I__1919 (
            .O(N__10786),
            .I(N__10783));
    LocalMux I__1918 (
            .O(N__10783),
            .I(beamY_RNIGO5PPVZ0Z_0));
    InMux I__1917 (
            .O(N__10780),
            .I(N__10777));
    LocalMux I__1916 (
            .O(N__10777),
            .I(N_345_0_0_1));
    CascadeMux I__1915 (
            .O(N__10774),
            .I(font_un28_pixel_29_cascade_));
    CascadeMux I__1914 (
            .O(N__10771),
            .I(un116_pixel_5_am_6_cascade_));
    InMux I__1913 (
            .O(N__10768),
            .I(N__10765));
    LocalMux I__1912 (
            .O(N__10765),
            .I(g1_1));
    CascadeMux I__1911 (
            .O(N__10762),
            .I(N__10759));
    InMux I__1910 (
            .O(N__10759),
            .I(N__10756));
    LocalMux I__1909 (
            .O(N__10756),
            .I(g0_0_x2_1));
    CascadeMux I__1908 (
            .O(N__10753),
            .I(un114_pixel_1_0_3__un116_pixel_2_ns_1Z0Z_2_cascade_));
    CascadeMux I__1907 (
            .O(N__10750),
            .I(un114_pixel_1_0_3__un116_pixel_5_ns_1Z0Z_2_cascade_));
    CascadeMux I__1906 (
            .O(N__10747),
            .I(N__10743));
    InMux I__1905 (
            .O(N__10746),
            .I(N__10739));
    InMux I__1904 (
            .O(N__10743),
            .I(N__10736));
    InMux I__1903 (
            .O(N__10742),
            .I(N__10732));
    LocalMux I__1902 (
            .O(N__10739),
            .I(N__10729));
    LocalMux I__1901 (
            .O(N__10736),
            .I(N__10726));
    InMux I__1900 (
            .O(N__10735),
            .I(N__10723));
    LocalMux I__1899 (
            .O(N__10732),
            .I(beamXZ0Z_9));
    Odrv4 I__1898 (
            .O(N__10729),
            .I(beamXZ0Z_9));
    Odrv4 I__1897 (
            .O(N__10726),
            .I(beamXZ0Z_9));
    LocalMux I__1896 (
            .O(N__10723),
            .I(beamXZ0Z_9));
    InMux I__1895 (
            .O(N__10714),
            .I(un5_visiblex_cry_8));
    CascadeMux I__1894 (
            .O(N__10711),
            .I(un116_pixel_3_bm_2_cascade_));
    CascadeMux I__1893 (
            .O(N__10708),
            .I(N__10705));
    InMux I__1892 (
            .O(N__10705),
            .I(N__10702));
    LocalMux I__1891 (
            .O(N__10702),
            .I(un114_pixel_1_0_3__N_5_1_0));
    CascadeMux I__1890 (
            .O(N__10699),
            .I(un114_pixel_1_0_3__un116_pixel_4_ns_1_0_7_cascade_));
    InMux I__1889 (
            .O(N__10696),
            .I(N__10693));
    LocalMux I__1888 (
            .O(N__10693),
            .I(un114_pixel_1_0_3__g2_1Z0Z_0));
    CascadeMux I__1887 (
            .O(N__10690),
            .I(N__10687));
    InMux I__1886 (
            .O(N__10687),
            .I(N__10683));
    CascadeMux I__1885 (
            .O(N__10686),
            .I(N__10680));
    LocalMux I__1884 (
            .O(N__10683),
            .I(N__10677));
    InMux I__1883 (
            .O(N__10680),
            .I(N__10674));
    Odrv12 I__1882 (
            .O(N__10677),
            .I(beamY_RNIH9THADZ0Z_4));
    LocalMux I__1881 (
            .O(N__10674),
            .I(beamY_RNIH9THADZ0Z_4));
    InMux I__1880 (
            .O(N__10669),
            .I(N__10659));
    InMux I__1879 (
            .O(N__10668),
            .I(N__10655));
    InMux I__1878 (
            .O(N__10667),
            .I(N__10652));
    InMux I__1877 (
            .O(N__10666),
            .I(N__10649));
    InMux I__1876 (
            .O(N__10665),
            .I(N__10646));
    InMux I__1875 (
            .O(N__10664),
            .I(N__10643));
    InMux I__1874 (
            .O(N__10663),
            .I(N__10637));
    InMux I__1873 (
            .O(N__10662),
            .I(N__10634));
    LocalMux I__1872 (
            .O(N__10659),
            .I(N__10628));
    InMux I__1871 (
            .O(N__10658),
            .I(N__10625));
    LocalMux I__1870 (
            .O(N__10655),
            .I(N__10618));
    LocalMux I__1869 (
            .O(N__10652),
            .I(N__10618));
    LocalMux I__1868 (
            .O(N__10649),
            .I(N__10618));
    LocalMux I__1867 (
            .O(N__10646),
            .I(N__10613));
    LocalMux I__1866 (
            .O(N__10643),
            .I(N__10613));
    InMux I__1865 (
            .O(N__10642),
            .I(N__10610));
    InMux I__1864 (
            .O(N__10641),
            .I(N__10605));
    InMux I__1863 (
            .O(N__10640),
            .I(N__10605));
    LocalMux I__1862 (
            .O(N__10637),
            .I(N__10602));
    LocalMux I__1861 (
            .O(N__10634),
            .I(N__10599));
    InMux I__1860 (
            .O(N__10633),
            .I(N__10596));
    CascadeMux I__1859 (
            .O(N__10632),
            .I(N__10592));
    InMux I__1858 (
            .O(N__10631),
            .I(N__10589));
    Span12Mux_s4_v I__1857 (
            .O(N__10628),
            .I(N__10584));
    LocalMux I__1856 (
            .O(N__10625),
            .I(N__10584));
    Span4Mux_v I__1855 (
            .O(N__10618),
            .I(N__10575));
    Span4Mux_v I__1854 (
            .O(N__10613),
            .I(N__10575));
    LocalMux I__1853 (
            .O(N__10610),
            .I(N__10575));
    LocalMux I__1852 (
            .O(N__10605),
            .I(N__10575));
    Span4Mux_h I__1851 (
            .O(N__10602),
            .I(N__10568));
    Span4Mux_h I__1850 (
            .O(N__10599),
            .I(N__10568));
    LocalMux I__1849 (
            .O(N__10596),
            .I(N__10568));
    InMux I__1848 (
            .O(N__10595),
            .I(N__10563));
    InMux I__1847 (
            .O(N__10592),
            .I(N__10563));
    LocalMux I__1846 (
            .O(N__10589),
            .I(beamYZ0Z_3));
    Odrv12 I__1845 (
            .O(N__10584),
            .I(beamYZ0Z_3));
    Odrv4 I__1844 (
            .O(N__10575),
            .I(beamYZ0Z_3));
    Odrv4 I__1843 (
            .O(N__10568),
            .I(beamYZ0Z_3));
    LocalMux I__1842 (
            .O(N__10563),
            .I(beamYZ0Z_3));
    CascadeMux I__1841 (
            .O(N__10552),
            .I(N__10545));
    InMux I__1840 (
            .O(N__10551),
            .I(N__10542));
    InMux I__1839 (
            .O(N__10550),
            .I(N__10539));
    InMux I__1838 (
            .O(N__10549),
            .I(N__10534));
    InMux I__1837 (
            .O(N__10548),
            .I(N__10534));
    InMux I__1836 (
            .O(N__10545),
            .I(N__10531));
    LocalMux I__1835 (
            .O(N__10542),
            .I(beamXZ0Z_1));
    LocalMux I__1834 (
            .O(N__10539),
            .I(beamXZ0Z_1));
    LocalMux I__1833 (
            .O(N__10534),
            .I(beamXZ0Z_1));
    LocalMux I__1832 (
            .O(N__10531),
            .I(beamXZ0Z_1));
    InMux I__1831 (
            .O(N__10522),
            .I(un5_visiblex_cry_0));
    CascadeMux I__1830 (
            .O(N__10519),
            .I(N__10513));
    InMux I__1829 (
            .O(N__10518),
            .I(N__10510));
    InMux I__1828 (
            .O(N__10517),
            .I(N__10505));
    InMux I__1827 (
            .O(N__10516),
            .I(N__10505));
    InMux I__1826 (
            .O(N__10513),
            .I(N__10502));
    LocalMux I__1825 (
            .O(N__10510),
            .I(beamXZ0Z_2));
    LocalMux I__1824 (
            .O(N__10505),
            .I(beamXZ0Z_2));
    LocalMux I__1823 (
            .O(N__10502),
            .I(beamXZ0Z_2));
    InMux I__1822 (
            .O(N__10495),
            .I(un5_visiblex_cry_1));
    CascadeMux I__1821 (
            .O(N__10492),
            .I(N__10487));
    CascadeMux I__1820 (
            .O(N__10491),
            .I(N__10482));
    CascadeMux I__1819 (
            .O(N__10490),
            .I(N__10479));
    InMux I__1818 (
            .O(N__10487),
            .I(N__10476));
    InMux I__1817 (
            .O(N__10486),
            .I(N__10473));
    InMux I__1816 (
            .O(N__10485),
            .I(N__10468));
    InMux I__1815 (
            .O(N__10482),
            .I(N__10468));
    InMux I__1814 (
            .O(N__10479),
            .I(N__10465));
    LocalMux I__1813 (
            .O(N__10476),
            .I(beamXZ0Z_3));
    LocalMux I__1812 (
            .O(N__10473),
            .I(beamXZ0Z_3));
    LocalMux I__1811 (
            .O(N__10468),
            .I(beamXZ0Z_3));
    LocalMux I__1810 (
            .O(N__10465),
            .I(beamXZ0Z_3));
    InMux I__1809 (
            .O(N__10456),
            .I(un5_visiblex_cry_2));
    CascadeMux I__1808 (
            .O(N__10453),
            .I(N__10445));
    InMux I__1807 (
            .O(N__10452),
            .I(N__10442));
    InMux I__1806 (
            .O(N__10451),
            .I(N__10439));
    InMux I__1805 (
            .O(N__10450),
            .I(N__10436));
    InMux I__1804 (
            .O(N__10449),
            .I(N__10431));
    InMux I__1803 (
            .O(N__10448),
            .I(N__10431));
    InMux I__1802 (
            .O(N__10445),
            .I(N__10428));
    LocalMux I__1801 (
            .O(N__10442),
            .I(beamXZ0Z_4));
    LocalMux I__1800 (
            .O(N__10439),
            .I(beamXZ0Z_4));
    LocalMux I__1799 (
            .O(N__10436),
            .I(beamXZ0Z_4));
    LocalMux I__1798 (
            .O(N__10431),
            .I(beamXZ0Z_4));
    LocalMux I__1797 (
            .O(N__10428),
            .I(beamXZ0Z_4));
    InMux I__1796 (
            .O(N__10417),
            .I(un5_visiblex_cry_3));
    InMux I__1795 (
            .O(N__10414),
            .I(N__10407));
    InMux I__1794 (
            .O(N__10413),
            .I(N__10404));
    InMux I__1793 (
            .O(N__10412),
            .I(N__10401));
    CascadeMux I__1792 (
            .O(N__10411),
            .I(N__10398));
    CascadeMux I__1791 (
            .O(N__10410),
            .I(N__10394));
    LocalMux I__1790 (
            .O(N__10407),
            .I(N__10387));
    LocalMux I__1789 (
            .O(N__10404),
            .I(N__10387));
    LocalMux I__1788 (
            .O(N__10401),
            .I(N__10387));
    InMux I__1787 (
            .O(N__10398),
            .I(N__10382));
    InMux I__1786 (
            .O(N__10397),
            .I(N__10382));
    InMux I__1785 (
            .O(N__10394),
            .I(N__10379));
    Odrv4 I__1784 (
            .O(N__10387),
            .I(beamXZ0Z_5));
    LocalMux I__1783 (
            .O(N__10382),
            .I(beamXZ0Z_5));
    LocalMux I__1782 (
            .O(N__10379),
            .I(beamXZ0Z_5));
    InMux I__1781 (
            .O(N__10372),
            .I(un5_visiblex_cry_4));
    CascadeMux I__1780 (
            .O(N__10369),
            .I(N__10361));
    InMux I__1779 (
            .O(N__10368),
            .I(N__10358));
    InMux I__1778 (
            .O(N__10367),
            .I(N__10355));
    InMux I__1777 (
            .O(N__10366),
            .I(N__10352));
    InMux I__1776 (
            .O(N__10365),
            .I(N__10347));
    InMux I__1775 (
            .O(N__10364),
            .I(N__10347));
    InMux I__1774 (
            .O(N__10361),
            .I(N__10344));
    LocalMux I__1773 (
            .O(N__10358),
            .I(beamXZ0Z_6));
    LocalMux I__1772 (
            .O(N__10355),
            .I(beamXZ0Z_6));
    LocalMux I__1771 (
            .O(N__10352),
            .I(beamXZ0Z_6));
    LocalMux I__1770 (
            .O(N__10347),
            .I(beamXZ0Z_6));
    LocalMux I__1769 (
            .O(N__10344),
            .I(beamXZ0Z_6));
    InMux I__1768 (
            .O(N__10333),
            .I(un5_visiblex_cry_5));
    CascadeMux I__1767 (
            .O(N__10330),
            .I(N__10326));
    CascadeMux I__1766 (
            .O(N__10329),
            .I(N__10323));
    InMux I__1765 (
            .O(N__10326),
            .I(N__10316));
    InMux I__1764 (
            .O(N__10323),
            .I(N__10316));
    InMux I__1763 (
            .O(N__10322),
            .I(N__10313));
    InMux I__1762 (
            .O(N__10321),
            .I(N__10308));
    LocalMux I__1761 (
            .O(N__10316),
            .I(N__10305));
    LocalMux I__1760 (
            .O(N__10313),
            .I(N__10302));
    InMux I__1759 (
            .O(N__10312),
            .I(N__10299));
    InMux I__1758 (
            .O(N__10311),
            .I(N__10296));
    LocalMux I__1757 (
            .O(N__10308),
            .I(beamXZ0Z_7));
    Odrv4 I__1756 (
            .O(N__10305),
            .I(beamXZ0Z_7));
    Odrv4 I__1755 (
            .O(N__10302),
            .I(beamXZ0Z_7));
    LocalMux I__1754 (
            .O(N__10299),
            .I(beamXZ0Z_7));
    LocalMux I__1753 (
            .O(N__10296),
            .I(beamXZ0Z_7));
    InMux I__1752 (
            .O(N__10285),
            .I(un5_visiblex_cry_6));
    CascadeMux I__1751 (
            .O(N__10282),
            .I(N__10278));
    InMux I__1750 (
            .O(N__10281),
            .I(N__10274));
    InMux I__1749 (
            .O(N__10278),
            .I(N__10270));
    InMux I__1748 (
            .O(N__10277),
            .I(N__10267));
    LocalMux I__1747 (
            .O(N__10274),
            .I(N__10264));
    InMux I__1746 (
            .O(N__10273),
            .I(N__10261));
    LocalMux I__1745 (
            .O(N__10270),
            .I(N__10258));
    LocalMux I__1744 (
            .O(N__10267),
            .I(beamXZ0Z_8));
    Odrv4 I__1743 (
            .O(N__10264),
            .I(beamXZ0Z_8));
    LocalMux I__1742 (
            .O(N__10261),
            .I(beamXZ0Z_8));
    Odrv4 I__1741 (
            .O(N__10258),
            .I(beamXZ0Z_8));
    InMux I__1740 (
            .O(N__10249),
            .I(bfn_6_11_0_));
    InMux I__1739 (
            .O(N__10246),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_4));
    InMux I__1738 (
            .O(N__10243),
            .I(N__10240));
    LocalMux I__1737 (
            .O(N__10240),
            .I(un1_beamxlt10_0));
    CascadeMux I__1736 (
            .O(N__10237),
            .I(N__10232));
    InMux I__1735 (
            .O(N__10236),
            .I(N__10228));
    CascadeMux I__1734 (
            .O(N__10235),
            .I(N__10225));
    InMux I__1733 (
            .O(N__10232),
            .I(N__10222));
    InMux I__1732 (
            .O(N__10231),
            .I(N__10219));
    LocalMux I__1731 (
            .O(N__10228),
            .I(N__10216));
    InMux I__1730 (
            .O(N__10225),
            .I(N__10213));
    LocalMux I__1729 (
            .O(N__10222),
            .I(N__10210));
    LocalMux I__1728 (
            .O(N__10219),
            .I(beamXZ0Z_10));
    Odrv4 I__1727 (
            .O(N__10216),
            .I(beamXZ0Z_10));
    LocalMux I__1726 (
            .O(N__10213),
            .I(beamXZ0Z_10));
    Odrv4 I__1725 (
            .O(N__10210),
            .I(beamXZ0Z_10));
    CascadeMux I__1724 (
            .O(N__10201),
            .I(un114_pixel_1_0_3__un3_beamxZ0Z_5_cascade_));
    InMux I__1723 (
            .O(N__10198),
            .I(N__10195));
    LocalMux I__1722 (
            .O(N__10195),
            .I(N__10192));
    Odrv4 I__1721 (
            .O(N__10192),
            .I(un114_pixel_1_0_3__un3_beamxZ0Z_7));
    InMux I__1720 (
            .O(N__10189),
            .I(N__10183));
    InMux I__1719 (
            .O(N__10188),
            .I(N__10183));
    LocalMux I__1718 (
            .O(N__10183),
            .I(un18_beamylt4));
    InMux I__1717 (
            .O(N__10180),
            .I(N__10176));
    InMux I__1716 (
            .O(N__10179),
            .I(N__10171));
    LocalMux I__1715 (
            .O(N__10176),
            .I(N__10168));
    InMux I__1714 (
            .O(N__10175),
            .I(N__10163));
    InMux I__1713 (
            .O(N__10174),
            .I(N__10163));
    LocalMux I__1712 (
            .O(N__10171),
            .I(N__10160));
    Odrv4 I__1711 (
            .O(N__10168),
            .I(charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO));
    LocalMux I__1710 (
            .O(N__10163),
            .I(charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO));
    Odrv4 I__1709 (
            .O(N__10160),
            .I(charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO));
    CascadeMux I__1708 (
            .O(N__10153),
            .I(N__10150));
    InMux I__1707 (
            .O(N__10150),
            .I(N__10147));
    LocalMux I__1706 (
            .O(N__10147),
            .I(charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKFZ0));
    InMux I__1705 (
            .O(N__10144),
            .I(N__10141));
    LocalMux I__1704 (
            .O(N__10141),
            .I(charx_if_generate_plus_mult1_un19_sum_i));
    InMux I__1703 (
            .O(N__10138),
            .I(N__10131));
    InMux I__1702 (
            .O(N__10137),
            .I(N__10128));
    InMux I__1701 (
            .O(N__10136),
            .I(N__10125));
    InMux I__1700 (
            .O(N__10135),
            .I(N__10120));
    InMux I__1699 (
            .O(N__10134),
            .I(N__10120));
    LocalMux I__1698 (
            .O(N__10131),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    LocalMux I__1697 (
            .O(N__10128),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    LocalMux I__1696 (
            .O(N__10125),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    LocalMux I__1695 (
            .O(N__10120),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1));
    CascadeMux I__1694 (
            .O(N__10111),
            .I(N__10106));
    InMux I__1693 (
            .O(N__10110),
            .I(N__10103));
    InMux I__1692 (
            .O(N__10109),
            .I(N__10098));
    InMux I__1691 (
            .O(N__10106),
            .I(N__10098));
    LocalMux I__1690 (
            .O(N__10103),
            .I(beamY_RNI2MTA1Z0Z_9));
    LocalMux I__1689 (
            .O(N__10098),
            .I(beamY_RNI2MTA1Z0Z_9));
    CascadeMux I__1688 (
            .O(N__10093),
            .I(chary_if_generate_plus_mult1_un54_sum_c4_cascade_));
    InMux I__1687 (
            .O(N__10090),
            .I(N__10072));
    InMux I__1686 (
            .O(N__10089),
            .I(N__10072));
    InMux I__1685 (
            .O(N__10088),
            .I(N__10072));
    InMux I__1684 (
            .O(N__10087),
            .I(N__10072));
    InMux I__1683 (
            .O(N__10086),
            .I(N__10065));
    InMux I__1682 (
            .O(N__10085),
            .I(N__10065));
    InMux I__1681 (
            .O(N__10084),
            .I(N__10065));
    InMux I__1680 (
            .O(N__10083),
            .I(N__10060));
    InMux I__1679 (
            .O(N__10082),
            .I(N__10060));
    InMux I__1678 (
            .O(N__10081),
            .I(N__10057));
    LocalMux I__1677 (
            .O(N__10072),
            .I(beamY_RNICG8P9Z0Z_7));
    LocalMux I__1676 (
            .O(N__10065),
            .I(beamY_RNICG8P9Z0Z_7));
    LocalMux I__1675 (
            .O(N__10060),
            .I(beamY_RNICG8P9Z0Z_7));
    LocalMux I__1674 (
            .O(N__10057),
            .I(beamY_RNICG8P9Z0Z_7));
    InMux I__1673 (
            .O(N__10048),
            .I(N__10036));
    InMux I__1672 (
            .O(N__10047),
            .I(N__10036));
    InMux I__1671 (
            .O(N__10046),
            .I(N__10036));
    InMux I__1670 (
            .O(N__10045),
            .I(N__10031));
    InMux I__1669 (
            .O(N__10044),
            .I(N__10026));
    InMux I__1668 (
            .O(N__10043),
            .I(N__10026));
    LocalMux I__1667 (
            .O(N__10036),
            .I(N__10023));
    InMux I__1666 (
            .O(N__10035),
            .I(N__10018));
    InMux I__1665 (
            .O(N__10034),
            .I(N__10018));
    LocalMux I__1664 (
            .O(N__10031),
            .I(N__10013));
    LocalMux I__1663 (
            .O(N__10026),
            .I(N__10013));
    Span4Mux_h I__1662 (
            .O(N__10023),
            .I(N__10010));
    LocalMux I__1661 (
            .O(N__10018),
            .I(N__10005));
    Span4Mux_s2_v I__1660 (
            .O(N__10013),
            .I(N__10005));
    Odrv4 I__1659 (
            .O(N__10010),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    Odrv4 I__1658 (
            .O(N__10005),
            .I(chary_if_generate_plus_mult1_un61_sum_axbxc5_1));
    CascadeMux I__1657 (
            .O(N__10000),
            .I(un3_beamx_0_cascade_));
    InMux I__1656 (
            .O(N__9997),
            .I(N__9991));
    InMux I__1655 (
            .O(N__9996),
            .I(N__9991));
    LocalMux I__1654 (
            .O(N__9991),
            .I(un1_beamx_2));
    IoInMux I__1653 (
            .O(N__9988),
            .I(N__9985));
    LocalMux I__1652 (
            .O(N__9985),
            .I(N__9982));
    Span4Mux_s2_v I__1651 (
            .O(N__9982),
            .I(N__9979));
    Span4Mux_v I__1650 (
            .O(N__9979),
            .I(N__9976));
    Odrv4 I__1649 (
            .O(N__9976),
            .I(HSync_c));
    InMux I__1648 (
            .O(N__9973),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_1));
    InMux I__1647 (
            .O(N__9970),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_2));
    CascadeMux I__1646 (
            .O(N__9967),
            .I(N__9964));
    InMux I__1645 (
            .O(N__9964),
            .I(N__9961));
    LocalMux I__1644 (
            .O(N__9961),
            .I(N__9958));
    Odrv4 I__1643 (
            .O(N__9958),
            .I(charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8VZ0));
    InMux I__1642 (
            .O(N__9955),
            .I(charx_if_generate_plus_mult1_un26_sum_cry_3));
    CascadeMux I__1641 (
            .O(N__9952),
            .I(N__9949));
    InMux I__1640 (
            .O(N__9949),
            .I(N__9946));
    LocalMux I__1639 (
            .O(N__9946),
            .I(g0_3_2));
    CascadeMux I__1638 (
            .O(N__9943),
            .I(beamY_RNIARUFBZ0Z_5_cascade_));
    InMux I__1637 (
            .O(N__9940),
            .I(N__9937));
    LocalMux I__1636 (
            .O(N__9937),
            .I(beamY_RNIGS0LBZ0Z_5));
    InMux I__1635 (
            .O(N__9934),
            .I(N__9928));
    InMux I__1634 (
            .O(N__9933),
            .I(N__9925));
    InMux I__1633 (
            .O(N__9932),
            .I(N__9920));
    CascadeMux I__1632 (
            .O(N__9931),
            .I(N__9917));
    LocalMux I__1631 (
            .O(N__9928),
            .I(N__9912));
    LocalMux I__1630 (
            .O(N__9925),
            .I(N__9912));
    InMux I__1629 (
            .O(N__9924),
            .I(N__9903));
    InMux I__1628 (
            .O(N__9923),
            .I(N__9900));
    LocalMux I__1627 (
            .O(N__9920),
            .I(N__9897));
    InMux I__1626 (
            .O(N__9917),
            .I(N__9894));
    Span4Mux_h I__1625 (
            .O(N__9912),
            .I(N__9891));
    InMux I__1624 (
            .O(N__9911),
            .I(N__9882));
    InMux I__1623 (
            .O(N__9910),
            .I(N__9882));
    InMux I__1622 (
            .O(N__9909),
            .I(N__9882));
    InMux I__1621 (
            .O(N__9908),
            .I(N__9882));
    InMux I__1620 (
            .O(N__9907),
            .I(N__9877));
    InMux I__1619 (
            .O(N__9906),
            .I(N__9877));
    LocalMux I__1618 (
            .O(N__9903),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    LocalMux I__1617 (
            .O(N__9900),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    Odrv4 I__1616 (
            .O(N__9897),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    LocalMux I__1615 (
            .O(N__9894),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    Odrv4 I__1614 (
            .O(N__9891),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    LocalMux I__1613 (
            .O(N__9882),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    LocalMux I__1612 (
            .O(N__9877),
            .I(chary_if_generate_plus_mult1_un54_sum_c5));
    CascadeMux I__1611 (
            .O(N__9862),
            .I(chary_if_generate_plus_mult1_un54_sum_c5_cascade_));
    InMux I__1610 (
            .O(N__9859),
            .I(N__9852));
    InMux I__1609 (
            .O(N__9858),
            .I(N__9847));
    InMux I__1608 (
            .O(N__9857),
            .I(N__9847));
    InMux I__1607 (
            .O(N__9856),
            .I(N__9840));
    InMux I__1606 (
            .O(N__9855),
            .I(N__9840));
    LocalMux I__1605 (
            .O(N__9852),
            .I(N__9835));
    LocalMux I__1604 (
            .O(N__9847),
            .I(N__9835));
    InMux I__1603 (
            .O(N__9846),
            .I(N__9830));
    InMux I__1602 (
            .O(N__9845),
            .I(N__9830));
    LocalMux I__1601 (
            .O(N__9840),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0));
    Odrv4 I__1600 (
            .O(N__9835),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0));
    LocalMux I__1599 (
            .O(N__9830),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0));
    InMux I__1598 (
            .O(N__9823),
            .I(N__9820));
    LocalMux I__1597 (
            .O(N__9820),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0_0));
    InMux I__1596 (
            .O(N__9817),
            .I(N__9812));
    CascadeMux I__1595 (
            .O(N__9816),
            .I(N__9809));
    CascadeMux I__1594 (
            .O(N__9815),
            .I(N__9805));
    LocalMux I__1593 (
            .O(N__9812),
            .I(N__9800));
    InMux I__1592 (
            .O(N__9809),
            .I(N__9789));
    InMux I__1591 (
            .O(N__9808),
            .I(N__9789));
    InMux I__1590 (
            .O(N__9805),
            .I(N__9789));
    InMux I__1589 (
            .O(N__9804),
            .I(N__9789));
    InMux I__1588 (
            .O(N__9803),
            .I(N__9789));
    Odrv4 I__1587 (
            .O(N__9800),
            .I(beamY_RNIDO3IZ0Z_9));
    LocalMux I__1586 (
            .O(N__9789),
            .I(beamY_RNIDO3IZ0Z_9));
    InMux I__1585 (
            .O(N__9784),
            .I(N__9777));
    CascadeMux I__1584 (
            .O(N__9783),
            .I(N__9774));
    CascadeMux I__1583 (
            .O(N__9782),
            .I(N__9771));
    CascadeMux I__1582 (
            .O(N__9781),
            .I(N__9766));
    InMux I__1581 (
            .O(N__9780),
            .I(N__9757));
    LocalMux I__1580 (
            .O(N__9777),
            .I(N__9754));
    InMux I__1579 (
            .O(N__9774),
            .I(N__9751));
    InMux I__1578 (
            .O(N__9771),
            .I(N__9746));
    InMux I__1577 (
            .O(N__9770),
            .I(N__9746));
    InMux I__1576 (
            .O(N__9769),
            .I(N__9743));
    InMux I__1575 (
            .O(N__9766),
            .I(N__9740));
    InMux I__1574 (
            .O(N__9765),
            .I(N__9735));
    InMux I__1573 (
            .O(N__9764),
            .I(N__9730));
    InMux I__1572 (
            .O(N__9763),
            .I(N__9730));
    InMux I__1571 (
            .O(N__9762),
            .I(N__9725));
    InMux I__1570 (
            .O(N__9761),
            .I(N__9725));
    CascadeMux I__1569 (
            .O(N__9760),
            .I(N__9722));
    LocalMux I__1568 (
            .O(N__9757),
            .I(N__9715));
    Span4Mux_v I__1567 (
            .O(N__9754),
            .I(N__9715));
    LocalMux I__1566 (
            .O(N__9751),
            .I(N__9706));
    LocalMux I__1565 (
            .O(N__9746),
            .I(N__9706));
    LocalMux I__1564 (
            .O(N__9743),
            .I(N__9706));
    LocalMux I__1563 (
            .O(N__9740),
            .I(N__9706));
    CascadeMux I__1562 (
            .O(N__9739),
            .I(N__9703));
    CascadeMux I__1561 (
            .O(N__9738),
            .I(N__9700));
    LocalMux I__1560 (
            .O(N__9735),
            .I(N__9695));
    LocalMux I__1559 (
            .O(N__9730),
            .I(N__9690));
    LocalMux I__1558 (
            .O(N__9725),
            .I(N__9690));
    InMux I__1557 (
            .O(N__9722),
            .I(N__9685));
    InMux I__1556 (
            .O(N__9721),
            .I(N__9685));
    InMux I__1555 (
            .O(N__9720),
            .I(N__9682));
    Span4Mux_v I__1554 (
            .O(N__9715),
            .I(N__9677));
    Span4Mux_v I__1553 (
            .O(N__9706),
            .I(N__9677));
    InMux I__1552 (
            .O(N__9703),
            .I(N__9672));
    InMux I__1551 (
            .O(N__9700),
            .I(N__9672));
    InMux I__1550 (
            .O(N__9699),
            .I(N__9669));
    InMux I__1549 (
            .O(N__9698),
            .I(N__9666));
    Span4Mux_v I__1548 (
            .O(N__9695),
            .I(N__9661));
    Span4Mux_v I__1547 (
            .O(N__9690),
            .I(N__9661));
    LocalMux I__1546 (
            .O(N__9685),
            .I(N__9652));
    LocalMux I__1545 (
            .O(N__9682),
            .I(N__9652));
    Sp12to4 I__1544 (
            .O(N__9677),
            .I(N__9652));
    LocalMux I__1543 (
            .O(N__9672),
            .I(N__9652));
    LocalMux I__1542 (
            .O(N__9669),
            .I(N__9647));
    LocalMux I__1541 (
            .O(N__9666),
            .I(N__9647));
    Odrv4 I__1540 (
            .O(N__9661),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv12 I__1539 (
            .O(N__9652),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    Odrv12 I__1538 (
            .O(N__9647),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum));
    CascadeMux I__1537 (
            .O(N__9640),
            .I(N__9635));
    CascadeMux I__1536 (
            .O(N__9639),
            .I(N__9631));
    CascadeMux I__1535 (
            .O(N__9638),
            .I(N__9627));
    InMux I__1534 (
            .O(N__9635),
            .I(N__9621));
    InMux I__1533 (
            .O(N__9634),
            .I(N__9621));
    InMux I__1532 (
            .O(N__9631),
            .I(N__9618));
    InMux I__1531 (
            .O(N__9630),
            .I(N__9611));
    InMux I__1530 (
            .O(N__9627),
            .I(N__9611));
    InMux I__1529 (
            .O(N__9626),
            .I(N__9611));
    LocalMux I__1528 (
            .O(N__9621),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0));
    LocalMux I__1527 (
            .O(N__9618),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0));
    LocalMux I__1526 (
            .O(N__9611),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0));
    CascadeMux I__1525 (
            .O(N__9604),
            .I(N__9601));
    InMux I__1524 (
            .O(N__9601),
            .I(N__9598));
    LocalMux I__1523 (
            .O(N__9598),
            .I(N__9595));
    Odrv4 I__1522 (
            .O(N__9595),
            .I(g0_4_2));
    InMux I__1521 (
            .O(N__9592),
            .I(N__9584));
    InMux I__1520 (
            .O(N__9591),
            .I(N__9579));
    InMux I__1519 (
            .O(N__9590),
            .I(N__9579));
    InMux I__1518 (
            .O(N__9589),
            .I(N__9572));
    InMux I__1517 (
            .O(N__9588),
            .I(N__9572));
    InMux I__1516 (
            .O(N__9587),
            .I(N__9572));
    LocalMux I__1515 (
            .O(N__9584),
            .I(N__9565));
    LocalMux I__1514 (
            .O(N__9579),
            .I(N__9565));
    LocalMux I__1513 (
            .O(N__9572),
            .I(N__9562));
    InMux I__1512 (
            .O(N__9571),
            .I(N__9559));
    InMux I__1511 (
            .O(N__9570),
            .I(N__9556));
    Span4Mux_v I__1510 (
            .O(N__9565),
            .I(N__9551));
    Span4Mux_h I__1509 (
            .O(N__9562),
            .I(N__9551));
    LocalMux I__1508 (
            .O(N__9559),
            .I(N__9546));
    LocalMux I__1507 (
            .O(N__9556),
            .I(N__9546));
    Span4Mux_h I__1506 (
            .O(N__9551),
            .I(N__9530));
    Span4Mux_h I__1505 (
            .O(N__9546),
            .I(N__9530));
    InMux I__1504 (
            .O(N__9545),
            .I(N__9521));
    InMux I__1503 (
            .O(N__9544),
            .I(N__9521));
    InMux I__1502 (
            .O(N__9543),
            .I(N__9521));
    InMux I__1501 (
            .O(N__9542),
            .I(N__9521));
    InMux I__1500 (
            .O(N__9541),
            .I(N__9512));
    InMux I__1499 (
            .O(N__9540),
            .I(N__9512));
    InMux I__1498 (
            .O(N__9539),
            .I(N__9512));
    InMux I__1497 (
            .O(N__9538),
            .I(N__9512));
    InMux I__1496 (
            .O(N__9537),
            .I(N__9507));
    InMux I__1495 (
            .O(N__9536),
            .I(N__9507));
    InMux I__1494 (
            .O(N__9535),
            .I(N__9504));
    Span4Mux_v I__1493 (
            .O(N__9530),
            .I(N__9501));
    LocalMux I__1492 (
            .O(N__9521),
            .I(N__9496));
    LocalMux I__1491 (
            .O(N__9512),
            .I(N__9496));
    LocalMux I__1490 (
            .O(N__9507),
            .I(N__9491));
    LocalMux I__1489 (
            .O(N__9504),
            .I(N__9491));
    Odrv4 I__1488 (
            .O(N__9501),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    Odrv12 I__1487 (
            .O(N__9496),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    Odrv12 I__1486 (
            .O(N__9491),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum));
    CascadeMux I__1485 (
            .O(N__9484),
            .I(N__9481));
    InMux I__1484 (
            .O(N__9481),
            .I(N__9475));
    InMux I__1483 (
            .O(N__9480),
            .I(N__9468));
    InMux I__1482 (
            .O(N__9479),
            .I(N__9468));
    InMux I__1481 (
            .O(N__9478),
            .I(N__9468));
    LocalMux I__1480 (
            .O(N__9475),
            .I(chary_if_generate_plus_mult1_un54_sum_axb3));
    LocalMux I__1479 (
            .O(N__9468),
            .I(chary_if_generate_plus_mult1_un54_sum_axb3));
    InMux I__1478 (
            .O(N__9463),
            .I(N__9455));
    CascadeMux I__1477 (
            .O(N__9462),
            .I(N__9452));
    CascadeMux I__1476 (
            .O(N__9461),
            .I(N__9442));
    CascadeMux I__1475 (
            .O(N__9460),
            .I(N__9439));
    InMux I__1474 (
            .O(N__9459),
            .I(N__9434));
    InMux I__1473 (
            .O(N__9458),
            .I(N__9434));
    LocalMux I__1472 (
            .O(N__9455),
            .I(N__9431));
    InMux I__1471 (
            .O(N__9452),
            .I(N__9428));
    InMux I__1470 (
            .O(N__9451),
            .I(N__9422));
    InMux I__1469 (
            .O(N__9450),
            .I(N__9422));
    InMux I__1468 (
            .O(N__9449),
            .I(N__9413));
    InMux I__1467 (
            .O(N__9448),
            .I(N__9413));
    InMux I__1466 (
            .O(N__9447),
            .I(N__9413));
    InMux I__1465 (
            .O(N__9446),
            .I(N__9413));
    InMux I__1464 (
            .O(N__9445),
            .I(N__9408));
    InMux I__1463 (
            .O(N__9442),
            .I(N__9408));
    InMux I__1462 (
            .O(N__9439),
            .I(N__9405));
    LocalMux I__1461 (
            .O(N__9434),
            .I(N__9400));
    Span4Mux_v I__1460 (
            .O(N__9431),
            .I(N__9395));
    LocalMux I__1459 (
            .O(N__9428),
            .I(N__9395));
    InMux I__1458 (
            .O(N__9427),
            .I(N__9392));
    LocalMux I__1457 (
            .O(N__9422),
            .I(N__9389));
    LocalMux I__1456 (
            .O(N__9413),
            .I(N__9382));
    LocalMux I__1455 (
            .O(N__9408),
            .I(N__9382));
    LocalMux I__1454 (
            .O(N__9405),
            .I(N__9382));
    InMux I__1453 (
            .O(N__9404),
            .I(N__9377));
    InMux I__1452 (
            .O(N__9403),
            .I(N__9377));
    Span4Mux_v I__1451 (
            .O(N__9400),
            .I(N__9372));
    Span4Mux_v I__1450 (
            .O(N__9395),
            .I(N__9372));
    LocalMux I__1449 (
            .O(N__9392),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1448 (
            .O(N__9389),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv12 I__1447 (
            .O(N__9382),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    LocalMux I__1446 (
            .O(N__9377),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    Odrv4 I__1445 (
            .O(N__9372),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum));
    InMux I__1444 (
            .O(N__9361),
            .I(N__9354));
    InMux I__1443 (
            .O(N__9360),
            .I(N__9349));
    InMux I__1442 (
            .O(N__9359),
            .I(N__9349));
    InMux I__1441 (
            .O(N__9358),
            .I(N__9345));
    InMux I__1440 (
            .O(N__9357),
            .I(N__9342));
    LocalMux I__1439 (
            .O(N__9354),
            .I(N__9337));
    LocalMux I__1438 (
            .O(N__9349),
            .I(N__9337));
    InMux I__1437 (
            .O(N__9348),
            .I(N__9334));
    LocalMux I__1436 (
            .O(N__9345),
            .I(beamY_RNITFRN03Z0Z_5));
    LocalMux I__1435 (
            .O(N__9342),
            .I(beamY_RNITFRN03Z0Z_5));
    Odrv4 I__1434 (
            .O(N__9337),
            .I(beamY_RNITFRN03Z0Z_5));
    LocalMux I__1433 (
            .O(N__9334),
            .I(beamY_RNITFRN03Z0Z_5));
    InMux I__1432 (
            .O(N__9325),
            .I(N__9319));
    InMux I__1431 (
            .O(N__9324),
            .I(N__9314));
    InMux I__1430 (
            .O(N__9323),
            .I(N__9314));
    InMux I__1429 (
            .O(N__9322),
            .I(N__9311));
    LocalMux I__1428 (
            .O(N__9319),
            .I(N__9308));
    LocalMux I__1427 (
            .O(N__9314),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    LocalMux I__1426 (
            .O(N__9311),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    Odrv4 I__1425 (
            .O(N__9308),
            .I(chary_if_generate_plus_mult1_un75_sum_c5));
    CascadeMux I__1424 (
            .O(N__9301),
            .I(beamY_RNIH9THADZ0Z_4_cascade_));
    InMux I__1423 (
            .O(N__9298),
            .I(N__9292));
    CascadeMux I__1422 (
            .O(N__9297),
            .I(N__9289));
    InMux I__1421 (
            .O(N__9296),
            .I(N__9286));
    InMux I__1420 (
            .O(N__9295),
            .I(N__9283));
    LocalMux I__1419 (
            .O(N__9292),
            .I(N__9279));
    InMux I__1418 (
            .O(N__9289),
            .I(N__9276));
    LocalMux I__1417 (
            .O(N__9286),
            .I(N__9271));
    LocalMux I__1416 (
            .O(N__9283),
            .I(N__9271));
    InMux I__1415 (
            .O(N__9282),
            .I(N__9268));
    Odrv4 I__1414 (
            .O(N__9279),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0));
    LocalMux I__1413 (
            .O(N__9276),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0));
    Odrv4 I__1412 (
            .O(N__9271),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0));
    LocalMux I__1411 (
            .O(N__9268),
            .I(chary_if_generate_plus_mult1_un61_sum_axb3_0));
    InMux I__1410 (
            .O(N__9259),
            .I(N__9251));
    InMux I__1409 (
            .O(N__9258),
            .I(N__9248));
    InMux I__1408 (
            .O(N__9257),
            .I(N__9245));
    InMux I__1407 (
            .O(N__9256),
            .I(N__9240));
    InMux I__1406 (
            .O(N__9255),
            .I(N__9240));
    InMux I__1405 (
            .O(N__9254),
            .I(N__9237));
    LocalMux I__1404 (
            .O(N__9251),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d));
    LocalMux I__1403 (
            .O(N__9248),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d));
    LocalMux I__1402 (
            .O(N__9245),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d));
    LocalMux I__1401 (
            .O(N__9240),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d));
    LocalMux I__1400 (
            .O(N__9237),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d));
    CascadeMux I__1399 (
            .O(N__9226),
            .I(N__9223));
    InMux I__1398 (
            .O(N__9223),
            .I(N__9216));
    InMux I__1397 (
            .O(N__9222),
            .I(N__9216));
    InMux I__1396 (
            .O(N__9221),
            .I(N__9213));
    LocalMux I__1395 (
            .O(N__9216),
            .I(N__9210));
    LocalMux I__1394 (
            .O(N__9213),
            .I(N__9207));
    Span4Mux_v I__1393 (
            .O(N__9210),
            .I(N__9204));
    Odrv4 I__1392 (
            .O(N__9207),
            .I(beamY_RNIKHPCA1Z0Z_4));
    Odrv4 I__1391 (
            .O(N__9204),
            .I(beamY_RNIKHPCA1Z0Z_4));
    CascadeMux I__1390 (
            .O(N__9199),
            .I(chary_if_generate_plus_mult1_un61_sum_ac0_7_d_cascade_));
    InMux I__1389 (
            .O(N__9196),
            .I(N__9193));
    LocalMux I__1388 (
            .O(N__9193),
            .I(chary_if_generate_plus_mult1_un68_sum_axb4));
    InMux I__1387 (
            .O(N__9190),
            .I(N__9187));
    LocalMux I__1386 (
            .O(N__9187),
            .I(N__9181));
    InMux I__1385 (
            .O(N__9186),
            .I(N__9178));
    InMux I__1384 (
            .O(N__9185),
            .I(N__9173));
    InMux I__1383 (
            .O(N__9184),
            .I(N__9173));
    Span4Mux_v I__1382 (
            .O(N__9181),
            .I(N__9170));
    LocalMux I__1381 (
            .O(N__9178),
            .I(beamY_RNI2TEJF4Z0Z_4));
    LocalMux I__1380 (
            .O(N__9173),
            .I(beamY_RNI2TEJF4Z0Z_4));
    Odrv4 I__1379 (
            .O(N__9170),
            .I(beamY_RNI2TEJF4Z0Z_4));
    InMux I__1378 (
            .O(N__9163),
            .I(N__9154));
    InMux I__1377 (
            .O(N__9162),
            .I(N__9154));
    InMux I__1376 (
            .O(N__9161),
            .I(N__9151));
    InMux I__1375 (
            .O(N__9160),
            .I(N__9146));
    InMux I__1374 (
            .O(N__9159),
            .I(N__9146));
    LocalMux I__1373 (
            .O(N__9154),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    LocalMux I__1372 (
            .O(N__9151),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    LocalMux I__1371 (
            .O(N__9146),
            .I(chary_if_generate_plus_mult1_un68_sum_c4));
    InMux I__1370 (
            .O(N__9139),
            .I(N__9134));
    InMux I__1369 (
            .O(N__9138),
            .I(N__9131));
    InMux I__1368 (
            .O(N__9137),
            .I(N__9128));
    LocalMux I__1367 (
            .O(N__9134),
            .I(N__9125));
    LocalMux I__1366 (
            .O(N__9131),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_0));
    LocalMux I__1365 (
            .O(N__9128),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_0));
    Odrv4 I__1364 (
            .O(N__9125),
            .I(chary_if_generate_plus_mult1_un61_sum_axb4_0));
    CascadeMux I__1363 (
            .O(N__9118),
            .I(g0_0_x2_1_1_cascade_));
    CascadeMux I__1362 (
            .O(N__9115),
            .I(beamY_RNI2TEJF4Z0Z_4_cascade_));
    CascadeMux I__1361 (
            .O(N__9112),
            .I(N__9109));
    InMux I__1360 (
            .O(N__9109),
            .I(N__9106));
    LocalMux I__1359 (
            .O(N__9106),
            .I(un114_pixel_1_0_3__g0_8Z0Z_1));
    CascadeMux I__1358 (
            .O(N__9103),
            .I(chary_if_generate_plus_mult1_un61_sum_0_3_cascade_));
    CascadeMux I__1357 (
            .O(N__9100),
            .I(un114_pixel_1_0_3__g0_1Z0Z_1_cascade_));
    InMux I__1356 (
            .O(N__9097),
            .I(N__9094));
    LocalMux I__1355 (
            .O(N__9094),
            .I(chary_if_generate_plus_mult1_un61_sum_0_3));
    CascadeMux I__1354 (
            .O(N__9091),
            .I(un114_pixel_1_0_3__g0_3Z0Z_0_cascade_));
    InMux I__1353 (
            .O(N__9088),
            .I(N__9085));
    LocalMux I__1352 (
            .O(N__9085),
            .I(chary_if_generate_plus_mult1_un75_sum_i_0_5));
    InMux I__1351 (
            .O(N__9082),
            .I(N__9078));
    InMux I__1350 (
            .O(N__9081),
            .I(N__9075));
    LocalMux I__1349 (
            .O(N__9078),
            .I(chary_if_generate_plus_mult1_un68_sum_c4_0));
    LocalMux I__1348 (
            .O(N__9075),
            .I(chary_if_generate_plus_mult1_un68_sum_c4_0));
    CascadeMux I__1347 (
            .O(N__9070),
            .I(un114_pixel_1_0_3__g0Z0Z_1_cascade_));
    InMux I__1346 (
            .O(N__9067),
            .I(N__9064));
    LocalMux I__1345 (
            .O(N__9064),
            .I(chary_if_generate_plus_mult1_un68_sum_0_0_0_0_5));
    InMux I__1344 (
            .O(N__9061),
            .I(N__9058));
    LocalMux I__1343 (
            .O(N__9058),
            .I(g2));
    CascadeMux I__1342 (
            .O(N__9055),
            .I(un114_pixel_1_0_3__g0Z0Z_3_cascade_));
    CascadeMux I__1341 (
            .O(N__9052),
            .I(N__9049));
    InMux I__1340 (
            .O(N__9049),
            .I(N__9046));
    LocalMux I__1339 (
            .O(N__9046),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i));
    CascadeMux I__1338 (
            .O(N__9043),
            .I(N__9040));
    InMux I__1337 (
            .O(N__9040),
            .I(N__9037));
    LocalMux I__1336 (
            .O(N__9037),
            .I(N__9034));
    Odrv4 I__1335 (
            .O(N__9034),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i));
    InMux I__1334 (
            .O(N__9031),
            .I(N__9028));
    LocalMux I__1333 (
            .O(N__9028),
            .I(counter_27));
    InMux I__1332 (
            .O(N__9025),
            .I(N__9016));
    InMux I__1331 (
            .O(N__9024),
            .I(N__9016));
    InMux I__1330 (
            .O(N__9023),
            .I(N__9013));
    InMux I__1329 (
            .O(N__9022),
            .I(N__9008));
    InMux I__1328 (
            .O(N__9021),
            .I(N__9008));
    LocalMux I__1327 (
            .O(N__9016),
            .I(counterZ0Z_5));
    LocalMux I__1326 (
            .O(N__9013),
            .I(counterZ0Z_5));
    LocalMux I__1325 (
            .O(N__9008),
            .I(counterZ0Z_5));
    InMux I__1324 (
            .O(N__9001),
            .I(N__8995));
    InMux I__1323 (
            .O(N__9000),
            .I(N__8995));
    LocalMux I__1322 (
            .O(N__8995),
            .I(slaveselect_1_0_4));
    IoInMux I__1321 (
            .O(N__8992),
            .I(N__8988));
    IoInMux I__1320 (
            .O(N__8991),
            .I(N__8985));
    LocalMux I__1319 (
            .O(N__8988),
            .I(N__8980));
    LocalMux I__1318 (
            .O(N__8985),
            .I(N__8980));
    IoSpan4Mux I__1317 (
            .O(N__8980),
            .I(N__8977));
    Span4Mux_s3_v I__1316 (
            .O(N__8977),
            .I(N__8974));
    Odrv4 I__1315 (
            .O(N__8974),
            .I(un1_slaveselect_1_i));
    InMux I__1314 (
            .O(N__8971),
            .I(N__8959));
    InMux I__1313 (
            .O(N__8970),
            .I(N__8959));
    InMux I__1312 (
            .O(N__8969),
            .I(N__8959));
    InMux I__1311 (
            .O(N__8968),
            .I(N__8952));
    InMux I__1310 (
            .O(N__8967),
            .I(N__8952));
    InMux I__1309 (
            .O(N__8966),
            .I(N__8952));
    LocalMux I__1308 (
            .O(N__8959),
            .I(un3_slaveselect));
    LocalMux I__1307 (
            .O(N__8952),
            .I(un3_slaveselect));
    InMux I__1306 (
            .O(N__8947),
            .I(N__8944));
    LocalMux I__1305 (
            .O(N__8944),
            .I(counter_28));
    CascadeMux I__1304 (
            .O(N__8941),
            .I(N__8934));
    CascadeMux I__1303 (
            .O(N__8940),
            .I(N__8931));
    InMux I__1302 (
            .O(N__8939),
            .I(N__8928));
    InMux I__1301 (
            .O(N__8938),
            .I(N__8923));
    InMux I__1300 (
            .O(N__8937),
            .I(N__8923));
    InMux I__1299 (
            .O(N__8934),
            .I(N__8918));
    InMux I__1298 (
            .O(N__8931),
            .I(N__8918));
    LocalMux I__1297 (
            .O(N__8928),
            .I(counterZ0Z_4));
    LocalMux I__1296 (
            .O(N__8923),
            .I(counterZ0Z_4));
    LocalMux I__1295 (
            .O(N__8918),
            .I(counterZ0Z_4));
    CascadeMux I__1294 (
            .O(N__8911),
            .I(N__8904));
    CascadeMux I__1293 (
            .O(N__8910),
            .I(N__8901));
    CascadeMux I__1292 (
            .O(N__8909),
            .I(N__8895));
    InMux I__1291 (
            .O(N__8908),
            .I(N__8890));
    InMux I__1290 (
            .O(N__8907),
            .I(N__8883));
    InMux I__1289 (
            .O(N__8904),
            .I(N__8883));
    InMux I__1288 (
            .O(N__8901),
            .I(N__8883));
    InMux I__1287 (
            .O(N__8900),
            .I(N__8880));
    InMux I__1286 (
            .O(N__8899),
            .I(N__8869));
    InMux I__1285 (
            .O(N__8898),
            .I(N__8869));
    InMux I__1284 (
            .O(N__8895),
            .I(N__8869));
    InMux I__1283 (
            .O(N__8894),
            .I(N__8869));
    InMux I__1282 (
            .O(N__8893),
            .I(N__8869));
    LocalMux I__1281 (
            .O(N__8890),
            .I(slaveselectZ0));
    LocalMux I__1280 (
            .O(N__8883),
            .I(slaveselectZ0));
    LocalMux I__1279 (
            .O(N__8880),
            .I(slaveselectZ0));
    LocalMux I__1278 (
            .O(N__8869),
            .I(slaveselectZ0));
    CascadeMux I__1277 (
            .O(N__8860),
            .I(N__8855));
    InMux I__1276 (
            .O(N__8859),
            .I(N__8847));
    InMux I__1275 (
            .O(N__8858),
            .I(N__8844));
    InMux I__1274 (
            .O(N__8855),
            .I(N__8839));
    InMux I__1273 (
            .O(N__8854),
            .I(N__8839));
    InMux I__1272 (
            .O(N__8853),
            .I(N__8836));
    InMux I__1271 (
            .O(N__8852),
            .I(N__8829));
    InMux I__1270 (
            .O(N__8851),
            .I(N__8829));
    InMux I__1269 (
            .O(N__8850),
            .I(N__8829));
    LocalMux I__1268 (
            .O(N__8847),
            .I(un1_counter_0));
    LocalMux I__1267 (
            .O(N__8844),
            .I(un1_counter_0));
    LocalMux I__1266 (
            .O(N__8839),
            .I(un1_counter_0));
    LocalMux I__1265 (
            .O(N__8836),
            .I(un1_counter_0));
    LocalMux I__1264 (
            .O(N__8829),
            .I(un1_counter_0));
    IoInMux I__1263 (
            .O(N__8818),
            .I(N__8814));
    IoInMux I__1262 (
            .O(N__8817),
            .I(N__8811));
    LocalMux I__1261 (
            .O(N__8814),
            .I(N__8806));
    LocalMux I__1260 (
            .O(N__8811),
            .I(N__8806));
    Span4Mux_s2_v I__1259 (
            .O(N__8806),
            .I(N__8803));
    Sp12to4 I__1258 (
            .O(N__8803),
            .I(N__8799));
    InMux I__1257 (
            .O(N__8802),
            .I(N__8796));
    Odrv12 I__1256 (
            .O(N__8799),
            .I(nCS1_c));
    LocalMux I__1255 (
            .O(N__8796),
            .I(nCS1_c));
    SRMux I__1254 (
            .O(N__8791),
            .I(N__8788));
    LocalMux I__1253 (
            .O(N__8788),
            .I(N__8785));
    Span4Mux_h I__1252 (
            .O(N__8785),
            .I(N__8782));
    Odrv4 I__1251 (
            .O(N__8782),
            .I(nCS1_0_sqmuxa));
    InMux I__1250 (
            .O(N__8779),
            .I(un8_beamx_cry_6));
    InMux I__1249 (
            .O(N__8776),
            .I(un8_beamx_cry_7));
    InMux I__1248 (
            .O(N__8773),
            .I(bfn_5_10_0_));
    InMux I__1247 (
            .O(N__8770),
            .I(un8_beamx_cry_9));
    CascadeMux I__1246 (
            .O(N__8767),
            .I(N__8764));
    InMux I__1245 (
            .O(N__8764),
            .I(N__8761));
    LocalMux I__1244 (
            .O(N__8761),
            .I(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0));
    InMux I__1243 (
            .O(N__8758),
            .I(charx_if_generate_plus_mult1_un19_sum_cry_2));
    InMux I__1242 (
            .O(N__8755),
            .I(N__8752));
    LocalMux I__1241 (
            .O(N__8752),
            .I(un13_beamylt7));
    CascadeMux I__1240 (
            .O(N__8749),
            .I(N__8745));
    InMux I__1239 (
            .O(N__8748),
            .I(N__8740));
    InMux I__1238 (
            .O(N__8745),
            .I(N__8740));
    LocalMux I__1237 (
            .O(N__8740),
            .I(if_generate_plus_mult1_un75_sum_axbxc5));
    InMux I__1236 (
            .O(N__8737),
            .I(N__8733));
    InMux I__1235 (
            .O(N__8736),
            .I(N__8730));
    LocalMux I__1234 (
            .O(N__8733),
            .I(if_generate_plus_mult1_un75_sum_axbxc3));
    LocalMux I__1233 (
            .O(N__8730),
            .I(if_generate_plus_mult1_un75_sum_axbxc3));
    CascadeMux I__1232 (
            .O(N__8725),
            .I(row_1_if_generate_plus_mult1_un82_sum_axb4_i_cascade_));
    InMux I__1231 (
            .O(N__8722),
            .I(N__8719));
    LocalMux I__1230 (
            .O(N__8719),
            .I(row_1_if_generate_plus_mult1_un82_sum_ac0_7_0Z0Z_1));
    InMux I__1229 (
            .O(N__8716),
            .I(un8_beamx_cry_1));
    InMux I__1228 (
            .O(N__8713),
            .I(un8_beamx_cry_2));
    InMux I__1227 (
            .O(N__8710),
            .I(un8_beamx_cry_3));
    InMux I__1226 (
            .O(N__8707),
            .I(un8_beamx_cry_4));
    InMux I__1225 (
            .O(N__8704),
            .I(un8_beamx_cry_5));
    InMux I__1224 (
            .O(N__8701),
            .I(N__8692));
    InMux I__1223 (
            .O(N__8700),
            .I(N__8692));
    InMux I__1222 (
            .O(N__8699),
            .I(N__8692));
    LocalMux I__1221 (
            .O(N__8692),
            .I(chary_if_generate_plus_mult1_un47_sum_c5));
    CascadeMux I__1220 (
            .O(N__8689),
            .I(beamY_RNITURI3_0Z0Z_7_cascade_));
    InMux I__1219 (
            .O(N__8686),
            .I(N__8683));
    LocalMux I__1218 (
            .O(N__8683),
            .I(beamY_RNITURI3Z0Z_7));
    InMux I__1217 (
            .O(N__8680),
            .I(N__8677));
    LocalMux I__1216 (
            .O(N__8677),
            .I(un4_beamy_0));
    InMux I__1215 (
            .O(N__8674),
            .I(N__8671));
    LocalMux I__1214 (
            .O(N__8671),
            .I(un8_beamy));
    InMux I__1213 (
            .O(N__8668),
            .I(N__8665));
    LocalMux I__1212 (
            .O(N__8665),
            .I(un114_pixel_1_0_3__un15_beamyZ0Z_2));
    CascadeMux I__1211 (
            .O(N__8662),
            .I(un1_beamx_2_cascade_));
    CascadeMux I__1210 (
            .O(N__8659),
            .I(N__8656));
    InMux I__1209 (
            .O(N__8656),
            .I(N__8653));
    LocalMux I__1208 (
            .O(N__8653),
            .I(N__8650));
    Odrv4 I__1207 (
            .O(N__8650),
            .I(un114_pixel_1_0_3__un5_beamxZ0Z_3));
    InMux I__1206 (
            .O(N__8647),
            .I(N__8638));
    InMux I__1205 (
            .O(N__8646),
            .I(N__8635));
    InMux I__1204 (
            .O(N__8645),
            .I(N__8630));
    InMux I__1203 (
            .O(N__8644),
            .I(N__8630));
    InMux I__1202 (
            .O(N__8643),
            .I(N__8626));
    InMux I__1201 (
            .O(N__8642),
            .I(N__8621));
    InMux I__1200 (
            .O(N__8641),
            .I(N__8621));
    LocalMux I__1199 (
            .O(N__8638),
            .I(N__8617));
    LocalMux I__1198 (
            .O(N__8635),
            .I(N__8612));
    LocalMux I__1197 (
            .O(N__8630),
            .I(N__8612));
    InMux I__1196 (
            .O(N__8629),
            .I(N__8609));
    LocalMux I__1195 (
            .O(N__8626),
            .I(N__8602));
    LocalMux I__1194 (
            .O(N__8621),
            .I(N__8602));
    InMux I__1193 (
            .O(N__8620),
            .I(N__8596));
    Span4Mux_v I__1192 (
            .O(N__8617),
            .I(N__8589));
    Span4Mux_v I__1191 (
            .O(N__8612),
            .I(N__8589));
    LocalMux I__1190 (
            .O(N__8609),
            .I(N__8589));
    InMux I__1189 (
            .O(N__8608),
            .I(N__8584));
    InMux I__1188 (
            .O(N__8607),
            .I(N__8584));
    Span4Mux_h I__1187 (
            .O(N__8602),
            .I(N__8581));
    InMux I__1186 (
            .O(N__8601),
            .I(N__8574));
    InMux I__1185 (
            .O(N__8600),
            .I(N__8574));
    InMux I__1184 (
            .O(N__8599),
            .I(N__8574));
    LocalMux I__1183 (
            .O(N__8596),
            .I(beamYZ0Z_4));
    Odrv4 I__1182 (
            .O(N__8589),
            .I(beamYZ0Z_4));
    LocalMux I__1181 (
            .O(N__8584),
            .I(beamYZ0Z_4));
    Odrv4 I__1180 (
            .O(N__8581),
            .I(beamYZ0Z_4));
    LocalMux I__1179 (
            .O(N__8574),
            .I(beamYZ0Z_4));
    InMux I__1178 (
            .O(N__8563),
            .I(N__8560));
    LocalMux I__1177 (
            .O(N__8560),
            .I(un114_pixel_1_0_3__g0_1Z0Z_3));
    CascadeMux I__1176 (
            .O(N__8557),
            .I(un114_pixel_1_0_3__un18_beamylto9Z0Z_2_cascade_));
    InMux I__1175 (
            .O(N__8554),
            .I(N__8551));
    LocalMux I__1174 (
            .O(N__8551),
            .I(un18_beamylt10_0));
    CascadeMux I__1173 (
            .O(N__8548),
            .I(N__8542));
    CascadeMux I__1172 (
            .O(N__8547),
            .I(N__8539));
    InMux I__1171 (
            .O(N__8546),
            .I(N__8536));
    InMux I__1170 (
            .O(N__8545),
            .I(N__8533));
    InMux I__1169 (
            .O(N__8542),
            .I(N__8530));
    InMux I__1168 (
            .O(N__8539),
            .I(N__8527));
    LocalMux I__1167 (
            .O(N__8536),
            .I(N__8524));
    LocalMux I__1166 (
            .O(N__8533),
            .I(N__8515));
    LocalMux I__1165 (
            .O(N__8530),
            .I(N__8515));
    LocalMux I__1164 (
            .O(N__8527),
            .I(N__8515));
    Span4Mux_h I__1163 (
            .O(N__8524),
            .I(N__8512));
    InMux I__1162 (
            .O(N__8523),
            .I(N__8509));
    InMux I__1161 (
            .O(N__8522),
            .I(N__8506));
    Span4Mux_h I__1160 (
            .O(N__8515),
            .I(N__8501));
    Span4Mux_v I__1159 (
            .O(N__8512),
            .I(N__8501));
    LocalMux I__1158 (
            .O(N__8509),
            .I(N__8498));
    LocalMux I__1157 (
            .O(N__8506),
            .I(N__8495));
    Odrv4 I__1156 (
            .O(N__8501),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    Odrv4 I__1155 (
            .O(N__8498),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    Odrv12 I__1154 (
            .O(N__8495),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum));
    CascadeMux I__1153 (
            .O(N__8488),
            .I(beamY_RNINITP61Z0Z_5_cascade_));
    InMux I__1152 (
            .O(N__8485),
            .I(N__8482));
    LocalMux I__1151 (
            .O(N__8482),
            .I(beamY_RNINITP61_1Z0Z_5));
    InMux I__1150 (
            .O(N__8479),
            .I(N__8473));
    InMux I__1149 (
            .O(N__8478),
            .I(N__8473));
    LocalMux I__1148 (
            .O(N__8473),
            .I(chary_if_generate_plus_mult1_un40_sum_axb3));
    CascadeMux I__1147 (
            .O(N__8470),
            .I(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0_cascade_));
    InMux I__1146 (
            .O(N__8467),
            .I(N__8464));
    LocalMux I__1145 (
            .O(N__8464),
            .I(chary_if_generate_plus_mult1_un47_sum_axbxc5_2));
    CascadeMux I__1144 (
            .O(N__8461),
            .I(chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_));
    InMux I__1143 (
            .O(N__8458),
            .I(N__8446));
    InMux I__1142 (
            .O(N__8457),
            .I(N__8446));
    InMux I__1141 (
            .O(N__8456),
            .I(N__8446));
    InMux I__1140 (
            .O(N__8455),
            .I(N__8446));
    LocalMux I__1139 (
            .O(N__8446),
            .I(chary_if_generate_plus_mult1_un40_sum_c4));
    InMux I__1138 (
            .O(N__8443),
            .I(N__8440));
    LocalMux I__1137 (
            .O(N__8440),
            .I(un5_visibley_0_29));
    CascadeMux I__1136 (
            .O(N__8437),
            .I(chary_if_generate_plus_mult1_un61_sum_c5_cascade_));
    InMux I__1135 (
            .O(N__8434),
            .I(N__8428));
    InMux I__1134 (
            .O(N__8433),
            .I(N__8428));
    LocalMux I__1133 (
            .O(N__8428),
            .I(chary_if_generate_plus_mult1_un61_sum_0_1_5));
    CascadeMux I__1132 (
            .O(N__8425),
            .I(chary_if_generate_plus_mult1_un68_sum_c4_0_cascade_));
    InMux I__1131 (
            .O(N__8422),
            .I(N__8419));
    LocalMux I__1130 (
            .O(N__8419),
            .I(g0_0_3));
    CascadeMux I__1129 (
            .O(N__8416),
            .I(g1_0_cascade_));
    InMux I__1128 (
            .O(N__8413),
            .I(N__8410));
    LocalMux I__1127 (
            .O(N__8410),
            .I(N__8407));
    Odrv4 I__1126 (
            .O(N__8407),
            .I(un4_beamylt6));
    CascadeMux I__1125 (
            .O(N__8404),
            .I(chary_if_generate_plus_mult1_un75_sum_c5_N_9_cascade_));
    InMux I__1124 (
            .O(N__8401),
            .I(N__8398));
    LocalMux I__1123 (
            .O(N__8398),
            .I(g0_1_2));
    CascadeMux I__1122 (
            .O(N__8395),
            .I(N__8392));
    InMux I__1121 (
            .O(N__8392),
            .I(N__8389));
    LocalMux I__1120 (
            .O(N__8389),
            .I(N__8386));
    Span4Mux_h I__1119 (
            .O(N__8386),
            .I(N__8383));
    Span4Mux_v I__1118 (
            .O(N__8383),
            .I(N__8380));
    Odrv4 I__1117 (
            .O(N__8380),
            .I(g0_2_0));
    CascadeMux I__1116 (
            .O(N__8377),
            .I(N__8374));
    InMux I__1115 (
            .O(N__8374),
            .I(N__8371));
    LocalMux I__1114 (
            .O(N__8371),
            .I(chary_if_generate_plus_mult1_un61_sum_1_0_1_0_3));
    InMux I__1113 (
            .O(N__8368),
            .I(N__8363));
    InMux I__1112 (
            .O(N__8367),
            .I(N__8360));
    InMux I__1111 (
            .O(N__8366),
            .I(N__8357));
    LocalMux I__1110 (
            .O(N__8363),
            .I(counterZ0Z_3));
    LocalMux I__1109 (
            .O(N__8360),
            .I(counterZ0Z_3));
    LocalMux I__1108 (
            .O(N__8357),
            .I(counterZ0Z_3));
    CascadeMux I__1107 (
            .O(N__8350),
            .I(N__8344));
    CascadeMux I__1106 (
            .O(N__8349),
            .I(N__8341));
    InMux I__1105 (
            .O(N__8348),
            .I(N__8336));
    InMux I__1104 (
            .O(N__8347),
            .I(N__8336));
    InMux I__1103 (
            .O(N__8344),
            .I(N__8333));
    InMux I__1102 (
            .O(N__8341),
            .I(N__8330));
    LocalMux I__1101 (
            .O(N__8336),
            .I(counterZ0Z_1));
    LocalMux I__1100 (
            .O(N__8333),
            .I(counterZ0Z_1));
    LocalMux I__1099 (
            .O(N__8330),
            .I(counterZ0Z_1));
    CascadeMux I__1098 (
            .O(N__8323),
            .I(un1_counterlto3_0_cascade_));
    InMux I__1097 (
            .O(N__8320),
            .I(N__8313));
    InMux I__1096 (
            .O(N__8319),
            .I(N__8313));
    InMux I__1095 (
            .O(N__8318),
            .I(N__8310));
    LocalMux I__1094 (
            .O(N__8313),
            .I(N__8307));
    LocalMux I__1093 (
            .O(N__8310),
            .I(counterZ0Z_2));
    Odrv4 I__1092 (
            .O(N__8307),
            .I(counterZ0Z_2));
    CascadeMux I__1091 (
            .O(N__8302),
            .I(g0_0_1_cascade_));
    InMux I__1090 (
            .O(N__8299),
            .I(N__8296));
    LocalMux I__1089 (
            .O(N__8296),
            .I(chary_if_generate_plus_mult1_un61_sum_c5));
    InMux I__1088 (
            .O(N__8293),
            .I(counter_cry_3));
    InMux I__1087 (
            .O(N__8290),
            .I(counter_cry_4));
    CascadeMux I__1086 (
            .O(N__8287),
            .I(slaveselect_1_0_4_cascade_));
    InMux I__1085 (
            .O(N__8284),
            .I(N__8281));
    LocalMux I__1084 (
            .O(N__8281),
            .I(counter_30));
    CascadeMux I__1083 (
            .O(N__8278),
            .I(un3_slaveselect_cascade_));
    InMux I__1082 (
            .O(N__8275),
            .I(N__8272));
    LocalMux I__1081 (
            .O(N__8272),
            .I(counter_29));
    CascadeMux I__1080 (
            .O(N__8269),
            .I(counter_31_cascade_));
    InMux I__1079 (
            .O(N__8266),
            .I(N__8258));
    InMux I__1078 (
            .O(N__8265),
            .I(N__8258));
    InMux I__1077 (
            .O(N__8264),
            .I(N__8253));
    InMux I__1076 (
            .O(N__8263),
            .I(N__8253));
    LocalMux I__1075 (
            .O(N__8258),
            .I(counterZ0Z_0));
    LocalMux I__1074 (
            .O(N__8253),
            .I(counterZ0Z_0));
    CascadeMux I__1073 (
            .O(N__8248),
            .I(N__8245));
    InMux I__1072 (
            .O(N__8245),
            .I(N__8242));
    LocalMux I__1071 (
            .O(N__8242),
            .I(N__8239));
    Odrv4 I__1070 (
            .O(N__8239),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KCZ0Z4));
    InMux I__1069 (
            .O(N__8236),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1068 (
            .O(N__8233),
            .I(N__8230));
    InMux I__1067 (
            .O(N__8230),
            .I(N__8227));
    LocalMux I__1066 (
            .O(N__8227),
            .I(N__8224));
    Odrv4 I__1065 (
            .O(N__8224),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGSZ0Z6));
    InMux I__1064 (
            .O(N__8221),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1063 (
            .O(N__8218),
            .I(N__8215));
    LocalMux I__1062 (
            .O(N__8215),
            .I(N__8212));
    Odrv4 I__1061 (
            .O(N__8212),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__1060 (
            .O(N__8209),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__1059 (
            .O(N__8206),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7));
    InMux I__1058 (
            .O(N__8203),
            .I(N__8196));
    InMux I__1057 (
            .O(N__8202),
            .I(N__8196));
    InMux I__1056 (
            .O(N__8201),
            .I(N__8193));
    LocalMux I__1055 (
            .O(N__8196),
            .I(N__8190));
    LocalMux I__1054 (
            .O(N__8193),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7));
    Odrv4 I__1053 (
            .O(N__8190),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7));
    InMux I__1052 (
            .O(N__8185),
            .I(N__8179));
    InMux I__1051 (
            .O(N__8184),
            .I(N__8179));
    LocalMux I__1050 (
            .O(N__8179),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8));
    InMux I__1049 (
            .O(N__8176),
            .I(counter_cry_1));
    InMux I__1048 (
            .O(N__8173),
            .I(counter_cry_2));
    CascadeMux I__1047 (
            .O(N__8170),
            .I(N__8167));
    InMux I__1046 (
            .O(N__8167),
            .I(N__8164));
    LocalMux I__1045 (
            .O(N__8164),
            .I(N__8161));
    Odrv12 I__1044 (
            .O(N__8161),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5_0_nsZ0Z_1));
    CascadeMux I__1043 (
            .O(N__8158),
            .I(N__8154));
    InMux I__1042 (
            .O(N__8157),
            .I(N__8149));
    InMux I__1041 (
            .O(N__8154),
            .I(N__8144));
    InMux I__1040 (
            .O(N__8153),
            .I(N__8144));
    InMux I__1039 (
            .O(N__8152),
            .I(N__8141));
    LocalMux I__1038 (
            .O(N__8149),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    LocalMux I__1037 (
            .O(N__8144),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    LocalMux I__1036 (
            .O(N__8141),
            .I(row_1_if_generate_plus_mult1_un68_sum_c5));
    CascadeMux I__1035 (
            .O(N__8134),
            .I(row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0_cascade_));
    InMux I__1034 (
            .O(N__8131),
            .I(N__8128));
    LocalMux I__1033 (
            .O(N__8128),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5));
    InMux I__1032 (
            .O(N__8125),
            .I(N__8121));
    InMux I__1031 (
            .O(N__8124),
            .I(N__8118));
    LocalMux I__1030 (
            .O(N__8121),
            .I(if_generate_plus_mult1_un54_sum_axbxc3));
    LocalMux I__1029 (
            .O(N__8118),
            .I(if_generate_plus_mult1_un54_sum_axbxc3));
    CascadeMux I__1028 (
            .O(N__8113),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5_cascade_));
    InMux I__1027 (
            .O(N__8110),
            .I(N__8107));
    LocalMux I__1026 (
            .O(N__8107),
            .I(row_1_if_generate_plus_mult1_un61_sum_c5));
    CascadeMux I__1025 (
            .O(N__8104),
            .I(row_1_if_generate_plus_mult1_un61_sum_c5_cascade_));
    InMux I__1024 (
            .O(N__8101),
            .I(N__8098));
    LocalMux I__1023 (
            .O(N__8098),
            .I(row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0));
    InMux I__1022 (
            .O(N__8095),
            .I(N__8092));
    LocalMux I__1021 (
            .O(N__8092),
            .I(if_generate_plus_mult1_un68_sum_c5_0_bm));
    InMux I__1020 (
            .O(N__8089),
            .I(N__8086));
    LocalMux I__1019 (
            .O(N__8086),
            .I(N__8083));
    Odrv4 I__1018 (
            .O(N__8083),
            .I(row_1_if_generate_plus_mult1_un61_sum_ac0_7_c));
    InMux I__1017 (
            .O(N__8080),
            .I(N__8074));
    InMux I__1016 (
            .O(N__8079),
            .I(N__8074));
    LocalMux I__1015 (
            .O(N__8074),
            .I(row_1_if_generate_plus_mult1_un75_sum_cZ0Z4));
    CascadeMux I__1014 (
            .O(N__8071),
            .I(row_1_if_generate_plus_mult1_un75_sum_cZ0Z4_cascade_));
    CascadeMux I__1013 (
            .O(N__8068),
            .I(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_));
    InMux I__1012 (
            .O(N__8065),
            .I(N__8056));
    InMux I__1011 (
            .O(N__8064),
            .I(N__8056));
    InMux I__1010 (
            .O(N__8063),
            .I(N__8056));
    LocalMux I__1009 (
            .O(N__8056),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1));
    CascadeMux I__1008 (
            .O(N__8053),
            .I(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_));
    InMux I__1007 (
            .O(N__8050),
            .I(N__8041));
    InMux I__1006 (
            .O(N__8049),
            .I(N__8041));
    InMux I__1005 (
            .O(N__8048),
            .I(N__8041));
    LocalMux I__1004 (
            .O(N__8041),
            .I(if_generate_plus_mult1_un68_sum_axbxc3));
    CascadeMux I__1003 (
            .O(N__8038),
            .I(N__8035));
    InMux I__1002 (
            .O(N__8035),
            .I(N__8032));
    LocalMux I__1001 (
            .O(N__8032),
            .I(un5_visibley_c5));
    CascadeMux I__1000 (
            .O(N__8029),
            .I(un5_visibley_c5_cascade_));
    CascadeMux I__999 (
            .O(N__8026),
            .I(un114_pixel_1_0_3__un5_beamxZ0Z_5_cascade_));
    CascadeMux I__998 (
            .O(N__8023),
            .I(un114_pixel_1_0_3__g0_1Z0Z_0_cascade_));
    CascadeMux I__997 (
            .O(N__8020),
            .I(N__8017));
    InMux I__996 (
            .O(N__8017),
            .I(N__8014));
    LocalMux I__995 (
            .O(N__8014),
            .I(N__8011));
    Odrv4 I__994 (
            .O(N__8011),
            .I(un4_beamylt8_0));
    CascadeMux I__993 (
            .O(N__8008),
            .I(N__8005));
    InMux I__992 (
            .O(N__8005),
            .I(N__8001));
    InMux I__991 (
            .O(N__8004),
            .I(N__7998));
    LocalMux I__990 (
            .O(N__8001),
            .I(N__7995));
    LocalMux I__989 (
            .O(N__7998),
            .I(N__7991));
    Span4Mux_h I__988 (
            .O(N__7995),
            .I(N__7988));
    InMux I__987 (
            .O(N__7994),
            .I(N__7985));
    Odrv4 I__986 (
            .O(N__7991),
            .I(un5_visibley_c2));
    Odrv4 I__985 (
            .O(N__7988),
            .I(un5_visibley_c2));
    LocalMux I__984 (
            .O(N__7985),
            .I(un5_visibley_c2));
    InMux I__983 (
            .O(N__7978),
            .I(N__7972));
    InMux I__982 (
            .O(N__7977),
            .I(N__7969));
    InMux I__981 (
            .O(N__7976),
            .I(N__7964));
    InMux I__980 (
            .O(N__7975),
            .I(N__7964));
    LocalMux I__979 (
            .O(N__7972),
            .I(N__7961));
    LocalMux I__978 (
            .O(N__7969),
            .I(N__7956));
    LocalMux I__977 (
            .O(N__7964),
            .I(N__7956));
    Span4Mux_h I__976 (
            .O(N__7961),
            .I(N__7952));
    Span4Mux_h I__975 (
            .O(N__7956),
            .I(N__7949));
    InMux I__974 (
            .O(N__7955),
            .I(N__7946));
    Odrv4 I__973 (
            .O(N__7952),
            .I(un1_beamy_4));
    Odrv4 I__972 (
            .O(N__7949),
            .I(un1_beamy_4));
    LocalMux I__971 (
            .O(N__7946),
            .I(un1_beamy_4));
    InMux I__970 (
            .O(N__7939),
            .I(N__7933));
    InMux I__969 (
            .O(N__7938),
            .I(N__7926));
    InMux I__968 (
            .O(N__7937),
            .I(N__7926));
    InMux I__967 (
            .O(N__7936),
            .I(N__7926));
    LocalMux I__966 (
            .O(N__7933),
            .I(N__7917));
    LocalMux I__965 (
            .O(N__7926),
            .I(N__7917));
    InMux I__964 (
            .O(N__7925),
            .I(N__7912));
    InMux I__963 (
            .O(N__7924),
            .I(N__7912));
    CascadeMux I__962 (
            .O(N__7923),
            .I(N__7907));
    InMux I__961 (
            .O(N__7922),
            .I(N__7903));
    Span4Mux_h I__960 (
            .O(N__7917),
            .I(N__7900));
    LocalMux I__959 (
            .O(N__7912),
            .I(N__7897));
    InMux I__958 (
            .O(N__7911),
            .I(N__7894));
    InMux I__957 (
            .O(N__7910),
            .I(N__7887));
    InMux I__956 (
            .O(N__7907),
            .I(N__7887));
    InMux I__955 (
            .O(N__7906),
            .I(N__7887));
    LocalMux I__954 (
            .O(N__7903),
            .I(beamYZ0Z_8));
    Odrv4 I__953 (
            .O(N__7900),
            .I(beamYZ0Z_8));
    Odrv12 I__952 (
            .O(N__7897),
            .I(beamYZ0Z_8));
    LocalMux I__951 (
            .O(N__7894),
            .I(beamYZ0Z_8));
    LocalMux I__950 (
            .O(N__7887),
            .I(beamYZ0Z_8));
    InMux I__949 (
            .O(N__7876),
            .I(N__7867));
    InMux I__948 (
            .O(N__7875),
            .I(N__7860));
    InMux I__947 (
            .O(N__7874),
            .I(N__7860));
    InMux I__946 (
            .O(N__7873),
            .I(N__7860));
    InMux I__945 (
            .O(N__7872),
            .I(N__7853));
    InMux I__944 (
            .O(N__7871),
            .I(N__7853));
    InMux I__943 (
            .O(N__7870),
            .I(N__7853));
    LocalMux I__942 (
            .O(N__7867),
            .I(N__7845));
    LocalMux I__941 (
            .O(N__7860),
            .I(N__7845));
    LocalMux I__940 (
            .O(N__7853),
            .I(N__7845));
    InMux I__939 (
            .O(N__7852),
            .I(N__7841));
    Span4Mux_v I__938 (
            .O(N__7845),
            .I(N__7838));
    InMux I__937 (
            .O(N__7844),
            .I(N__7835));
    LocalMux I__936 (
            .O(N__7841),
            .I(beamYZ0Z_9));
    Odrv4 I__935 (
            .O(N__7838),
            .I(beamYZ0Z_9));
    LocalMux I__934 (
            .O(N__7835),
            .I(beamYZ0Z_9));
    CascadeMux I__933 (
            .O(N__7828),
            .I(un114_pixel_1_0_3__un8_beamylto9Z0Z_1_cascade_));
    InMux I__932 (
            .O(N__7825),
            .I(N__7820));
    InMux I__931 (
            .O(N__7824),
            .I(N__7811));
    InMux I__930 (
            .O(N__7823),
            .I(N__7811));
    LocalMux I__929 (
            .O(N__7820),
            .I(N__7806));
    InMux I__928 (
            .O(N__7819),
            .I(N__7797));
    InMux I__927 (
            .O(N__7818),
            .I(N__7797));
    InMux I__926 (
            .O(N__7817),
            .I(N__7797));
    InMux I__925 (
            .O(N__7816),
            .I(N__7797));
    LocalMux I__924 (
            .O(N__7811),
            .I(N__7794));
    CascadeMux I__923 (
            .O(N__7810),
            .I(N__7791));
    InMux I__922 (
            .O(N__7809),
            .I(N__7788));
    Span4Mux_v I__921 (
            .O(N__7806),
            .I(N__7783));
    LocalMux I__920 (
            .O(N__7797),
            .I(N__7783));
    Span4Mux_h I__919 (
            .O(N__7794),
            .I(N__7780));
    InMux I__918 (
            .O(N__7791),
            .I(N__7777));
    LocalMux I__917 (
            .O(N__7788),
            .I(beamYZ0Z_7));
    Odrv4 I__916 (
            .O(N__7783),
            .I(beamYZ0Z_7));
    Odrv4 I__915 (
            .O(N__7780),
            .I(beamYZ0Z_7));
    LocalMux I__914 (
            .O(N__7777),
            .I(beamYZ0Z_7));
    CascadeMux I__913 (
            .O(N__7768),
            .I(un114_pixel_1_0_3__un1_beamylto9Z0Z_0_cascade_));
    CascadeMux I__912 (
            .O(N__7765),
            .I(un4_beamylt6_cascade_));
    InMux I__911 (
            .O(N__7762),
            .I(N__7759));
    LocalMux I__910 (
            .O(N__7759),
            .I(N__7755));
    InMux I__909 (
            .O(N__7758),
            .I(N__7752));
    Odrv4 I__908 (
            .O(N__7755),
            .I(un5_visibley_ac0_11_d));
    LocalMux I__907 (
            .O(N__7752),
            .I(un5_visibley_ac0_11_d));
    InMux I__906 (
            .O(N__7747),
            .I(N__7744));
    LocalMux I__905 (
            .O(N__7744),
            .I(N__7740));
    InMux I__904 (
            .O(N__7743),
            .I(N__7737));
    Span4Mux_v I__903 (
            .O(N__7740),
            .I(N__7734));
    LocalMux I__902 (
            .O(N__7737),
            .I(N__7731));
    Odrv4 I__901 (
            .O(N__7734),
            .I(un5_visibley_ac0_11_0_1));
    Odrv4 I__900 (
            .O(N__7731),
            .I(un5_visibley_ac0_11_0_1));
    CascadeMux I__899 (
            .O(N__7726),
            .I(N__7723));
    InMux I__898 (
            .O(N__7723),
            .I(N__7720));
    LocalMux I__897 (
            .O(N__7720),
            .I(un114_pixel_1_0_3__un1_beamylto9_3));
    CascadeMux I__896 (
            .O(N__7717),
            .I(N__7714));
    InMux I__895 (
            .O(N__7714),
            .I(N__7711));
    LocalMux I__894 (
            .O(N__7711),
            .I(N__7705));
    InMux I__893 (
            .O(N__7710),
            .I(N__7702));
    InMux I__892 (
            .O(N__7709),
            .I(N__7697));
    InMux I__891 (
            .O(N__7708),
            .I(N__7697));
    Odrv4 I__890 (
            .O(N__7705),
            .I(beamY_fastZ0Z_2));
    LocalMux I__889 (
            .O(N__7702),
            .I(beamY_fastZ0Z_2));
    LocalMux I__888 (
            .O(N__7697),
            .I(beamY_fastZ0Z_2));
    InMux I__887 (
            .O(N__7690),
            .I(N__7684));
    InMux I__886 (
            .O(N__7689),
            .I(N__7684));
    LocalMux I__885 (
            .O(N__7684),
            .I(N__7678));
    InMux I__884 (
            .O(N__7683),
            .I(N__7673));
    InMux I__883 (
            .O(N__7682),
            .I(N__7673));
    InMux I__882 (
            .O(N__7681),
            .I(N__7670));
    Span4Mux_v I__881 (
            .O(N__7678),
            .I(N__7665));
    LocalMux I__880 (
            .O(N__7673),
            .I(N__7665));
    LocalMux I__879 (
            .O(N__7670),
            .I(N__7659));
    Span4Mux_h I__878 (
            .O(N__7665),
            .I(N__7656));
    InMux I__877 (
            .O(N__7664),
            .I(N__7651));
    InMux I__876 (
            .O(N__7663),
            .I(N__7651));
    InMux I__875 (
            .O(N__7662),
            .I(N__7648));
    Odrv4 I__874 (
            .O(N__7659),
            .I(beamYZ0Z_5));
    Odrv4 I__873 (
            .O(N__7656),
            .I(beamYZ0Z_5));
    LocalMux I__872 (
            .O(N__7651),
            .I(beamYZ0Z_5));
    LocalMux I__871 (
            .O(N__7648),
            .I(beamYZ0Z_5));
    InMux I__870 (
            .O(N__7639),
            .I(N__7635));
    CascadeMux I__869 (
            .O(N__7638),
            .I(N__7630));
    LocalMux I__868 (
            .O(N__7635),
            .I(N__7627));
    InMux I__867 (
            .O(N__7634),
            .I(N__7624));
    InMux I__866 (
            .O(N__7633),
            .I(N__7619));
    InMux I__865 (
            .O(N__7630),
            .I(N__7619));
    Odrv12 I__864 (
            .O(N__7627),
            .I(beamY_fastZ0Z_3));
    LocalMux I__863 (
            .O(N__7624),
            .I(beamY_fastZ0Z_3));
    LocalMux I__862 (
            .O(N__7619),
            .I(beamY_fastZ0Z_3));
    CascadeMux I__861 (
            .O(N__7612),
            .I(beamY_fast_RNIM4P7Z0Z_2_cascade_));
    InMux I__860 (
            .O(N__7609),
            .I(N__7601));
    InMux I__859 (
            .O(N__7608),
            .I(N__7601));
    InMux I__858 (
            .O(N__7607),
            .I(N__7597));
    InMux I__857 (
            .O(N__7606),
            .I(N__7594));
    LocalMux I__856 (
            .O(N__7601),
            .I(N__7591));
    InMux I__855 (
            .O(N__7600),
            .I(N__7585));
    LocalMux I__854 (
            .O(N__7597),
            .I(N__7580));
    LocalMux I__853 (
            .O(N__7594),
            .I(N__7580));
    Span4Mux_h I__852 (
            .O(N__7591),
            .I(N__7577));
    InMux I__851 (
            .O(N__7590),
            .I(N__7574));
    InMux I__850 (
            .O(N__7589),
            .I(N__7569));
    InMux I__849 (
            .O(N__7588),
            .I(N__7569));
    LocalMux I__848 (
            .O(N__7585),
            .I(beamYZ0Z_6));
    Odrv4 I__847 (
            .O(N__7580),
            .I(beamYZ0Z_6));
    Odrv4 I__846 (
            .O(N__7577),
            .I(beamYZ0Z_6));
    LocalMux I__845 (
            .O(N__7574),
            .I(beamYZ0Z_6));
    LocalMux I__844 (
            .O(N__7569),
            .I(beamYZ0Z_6));
    InMux I__843 (
            .O(N__7558),
            .I(N__7555));
    LocalMux I__842 (
            .O(N__7555),
            .I(chessboardpixel_un174_pixel_0_1));
    InMux I__841 (
            .O(N__7552),
            .I(N__7549));
    LocalMux I__840 (
            .O(N__7549),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__839 (
            .O(N__7546),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__838 (
            .O(N__7543),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__837 (
            .O(N__7540),
            .I(N__7534));
    InMux I__836 (
            .O(N__7539),
            .I(N__7534));
    LocalMux I__835 (
            .O(N__7534),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__834 (
            .O(N__7531),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7));
    CascadeMux I__833 (
            .O(N__7528),
            .I(N__7525));
    InMux I__832 (
            .O(N__7525),
            .I(N__7522));
    LocalMux I__831 (
            .O(N__7522),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHFZ0));
    InMux I__830 (
            .O(N__7519),
            .I(N__7516));
    LocalMux I__829 (
            .O(N__7516),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJZ0Z5));
    InMux I__828 (
            .O(N__7513),
            .I(N__7509));
    InMux I__827 (
            .O(N__7512),
            .I(N__7506));
    LocalMux I__826 (
            .O(N__7509),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0));
    LocalMux I__825 (
            .O(N__7506),
            .I(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0));
    InMux I__824 (
            .O(N__7501),
            .I(N__7498));
    LocalMux I__823 (
            .O(N__7498),
            .I(un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1Z0Z_1));
    CascadeMux I__822 (
            .O(N__7495),
            .I(chessboardpixel_un200_pixel_0_1_cascade_));
    InMux I__821 (
            .O(N__7492),
            .I(N__7489));
    LocalMux I__820 (
            .O(N__7489),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5));
    CascadeMux I__819 (
            .O(N__7486),
            .I(N__7480));
    InMux I__818 (
            .O(N__7485),
            .I(N__7477));
    InMux I__817 (
            .O(N__7484),
            .I(N__7472));
    InMux I__816 (
            .O(N__7483),
            .I(N__7472));
    InMux I__815 (
            .O(N__7480),
            .I(N__7469));
    LocalMux I__814 (
            .O(N__7477),
            .I(beamY_i_2));
    LocalMux I__813 (
            .O(N__7472),
            .I(beamY_i_2));
    LocalMux I__812 (
            .O(N__7469),
            .I(beamY_i_2));
    InMux I__811 (
            .O(N__7462),
            .I(N__7456));
    InMux I__810 (
            .O(N__7461),
            .I(N__7456));
    LocalMux I__809 (
            .O(N__7456),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81BZ0));
    InMux I__808 (
            .O(N__7453),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__807 (
            .O(N__7450),
            .I(N__7447));
    InMux I__806 (
            .O(N__7447),
            .I(N__7444));
    LocalMux I__805 (
            .O(N__7444),
            .I(N__7441));
    Odrv4 I__804 (
            .O(N__7441),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEGZ0Z5));
    InMux I__803 (
            .O(N__7438),
            .I(N__7432));
    InMux I__802 (
            .O(N__7437),
            .I(N__7432));
    LocalMux I__801 (
            .O(N__7432),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODGZ0));
    InMux I__800 (
            .O(N__7429),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__799 (
            .O(N__7426),
            .I(N__7423));
    LocalMux I__798 (
            .O(N__7423),
            .I(N__7420));
    Odrv4 I__797 (
            .O(N__7420),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87VZ0Z68));
    InMux I__796 (
            .O(N__7417),
            .I(N__7414));
    LocalMux I__795 (
            .O(N__7414),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4JZ0));
    InMux I__794 (
            .O(N__7411),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__793 (
            .O(N__7408),
            .I(N__7405));
    InMux I__792 (
            .O(N__7405),
            .I(N__7402));
    LocalMux I__791 (
            .O(N__7402),
            .I(N__7399));
    Odrv4 I__790 (
            .O(N__7399),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05UZ0Z8));
    CascadeMux I__789 (
            .O(N__7396),
            .I(N__7392));
    CascadeMux I__788 (
            .O(N__7395),
            .I(N__7388));
    InMux I__787 (
            .O(N__7392),
            .I(N__7377));
    InMux I__786 (
            .O(N__7391),
            .I(N__7377));
    InMux I__785 (
            .O(N__7388),
            .I(N__7377));
    InMux I__784 (
            .O(N__7387),
            .I(N__7377));
    InMux I__783 (
            .O(N__7386),
            .I(N__7374));
    LocalMux I__782 (
            .O(N__7377),
            .I(N__7371));
    LocalMux I__781 (
            .O(N__7374),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0));
    Odrv4 I__780 (
            .O(N__7371),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0));
    InMux I__779 (
            .O(N__7366),
            .I(N__7363));
    LocalMux I__778 (
            .O(N__7363),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__777 (
            .O(N__7360),
            .I(N__7357));
    LocalMux I__776 (
            .O(N__7357),
            .I(N__7354));
    Odrv4 I__775 (
            .O(N__7354),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__774 (
            .O(N__7351),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__773 (
            .O(N__7348),
            .I(N__7339));
    InMux I__772 (
            .O(N__7347),
            .I(N__7339));
    InMux I__771 (
            .O(N__7346),
            .I(N__7339));
    LocalMux I__770 (
            .O(N__7339),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGKZ0));
    CascadeMux I__769 (
            .O(N__7336),
            .I(N__7333));
    InMux I__768 (
            .O(N__7333),
            .I(N__7326));
    InMux I__767 (
            .O(N__7332),
            .I(N__7326));
    InMux I__766 (
            .O(N__7331),
            .I(N__7323));
    LocalMux I__765 (
            .O(N__7326),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1));
    LocalMux I__764 (
            .O(N__7323),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1));
    InMux I__763 (
            .O(N__7318),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4));
    InMux I__762 (
            .O(N__7315),
            .I(N__7312));
    LocalMux I__761 (
            .O(N__7312),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO));
    InMux I__760 (
            .O(N__7309),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__759 (
            .O(N__7306),
            .I(N__7303));
    LocalMux I__758 (
            .O(N__7303),
            .I(beamY_RNIFJ0L_0Z0Z_8));
    InMux I__757 (
            .O(N__7300),
            .I(N__7297));
    LocalMux I__756 (
            .O(N__7297),
            .I(beamY_RNI19IJ_0Z0Z_9));
    CascadeMux I__755 (
            .O(N__7294),
            .I(N__7290));
    InMux I__754 (
            .O(N__7293),
            .I(N__7280));
    InMux I__753 (
            .O(N__7290),
            .I(N__7280));
    InMux I__752 (
            .O(N__7289),
            .I(N__7280));
    InMux I__751 (
            .O(N__7288),
            .I(N__7277));
    InMux I__750 (
            .O(N__7287),
            .I(N__7274));
    LocalMux I__749 (
            .O(N__7280),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9));
    LocalMux I__748 (
            .O(N__7277),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9));
    LocalMux I__747 (
            .O(N__7274),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9));
    InMux I__746 (
            .O(N__7267),
            .I(N__7264));
    LocalMux I__745 (
            .O(N__7264),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7));
    CascadeMux I__744 (
            .O(N__7261),
            .I(beamY_i_2_cascade_));
    CascadeMux I__743 (
            .O(N__7258),
            .I(un114_pixel_1_0_3__chessboardpixel_un200_pixellto4Z0Z_1_cascade_));
    CascadeMux I__742 (
            .O(N__7255),
            .I(chessboardpixel_un200_pixellt10_cascade_));
    InMux I__741 (
            .O(N__7252),
            .I(N__7249));
    LocalMux I__740 (
            .O(N__7249),
            .I(un5_visibley_c6_0_0_0));
    CascadeMux I__739 (
            .O(N__7246),
            .I(beamY_fast_RNI35GAZ0Z_2_cascade_));
    InMux I__738 (
            .O(N__7243),
            .I(N__7239));
    InMux I__737 (
            .O(N__7242),
            .I(N__7236));
    LocalMux I__736 (
            .O(N__7239),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    LocalMux I__735 (
            .O(N__7236),
            .I(un21_beamy_cry_2_c_RNICOZ0Z83));
    InMux I__734 (
            .O(N__7231),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2));
    InMux I__733 (
            .O(N__7228),
            .I(N__7225));
    LocalMux I__732 (
            .O(N__7225),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2LZ0));
    InMux I__731 (
            .O(N__7222),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__730 (
            .O(N__7219),
            .I(N__7216));
    LocalMux I__729 (
            .O(N__7216),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO));
    InMux I__728 (
            .O(N__7213),
            .I(N__7210));
    LocalMux I__727 (
            .O(N__7210),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RCZ0));
    InMux I__726 (
            .O(N__7207),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__725 (
            .O(N__7204),
            .I(N__7200));
    InMux I__724 (
            .O(N__7203),
            .I(N__7197));
    LocalMux I__723 (
            .O(N__7200),
            .I(un21_beamy_cry_6_c_RNIK4DZ0Z3));
    LocalMux I__722 (
            .O(N__7197),
            .I(un21_beamy_cry_6_c_RNIK4DZ0Z3));
    CascadeMux I__721 (
            .O(N__7192),
            .I(N__7188));
    InMux I__720 (
            .O(N__7191),
            .I(N__7183));
    InMux I__719 (
            .O(N__7188),
            .I(N__7183));
    LocalMux I__718 (
            .O(N__7183),
            .I(beamY_fastZ0Z_7));
    InMux I__717 (
            .O(N__7180),
            .I(N__7177));
    LocalMux I__716 (
            .O(N__7177),
            .I(beamY_fastZ0Z_5));
    InMux I__715 (
            .O(N__7174),
            .I(N__7170));
    InMux I__714 (
            .O(N__7173),
            .I(N__7167));
    LocalMux I__713 (
            .O(N__7170),
            .I(un21_beamy_cry_1_c_RNIALZ0Z73));
    LocalMux I__712 (
            .O(N__7167),
            .I(un21_beamy_cry_1_c_RNIALZ0Z73));
    InMux I__711 (
            .O(N__7162),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__710 (
            .O(N__7159),
            .I(N__7156));
    LocalMux I__709 (
            .O(N__7156),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CRZ0Z2));
    InMux I__708 (
            .O(N__7153),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__707 (
            .O(N__7150),
            .I(N__7147));
    InMux I__706 (
            .O(N__7147),
            .I(N__7144));
    LocalMux I__705 (
            .O(N__7144),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGIZ0Z3));
    InMux I__704 (
            .O(N__7141),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__703 (
            .O(N__7138),
            .I(N__7135));
    InMux I__702 (
            .O(N__7135),
            .I(N__7132));
    LocalMux I__701 (
            .O(N__7132),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJZ0Z6874));
    InMux I__700 (
            .O(N__7129),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__699 (
            .O(N__7126),
            .I(N__7123));
    LocalMux I__698 (
            .O(N__7123),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__697 (
            .O(N__7120),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    CascadeMux I__696 (
            .O(N__7117),
            .I(N__7114));
    InMux I__695 (
            .O(N__7114),
            .I(N__7111));
    LocalMux I__694 (
            .O(N__7111),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0));
    CascadeMux I__693 (
            .O(N__7108),
            .I(N__7103));
    InMux I__692 (
            .O(N__7107),
            .I(N__7098));
    InMux I__691 (
            .O(N__7106),
            .I(N__7089));
    InMux I__690 (
            .O(N__7103),
            .I(N__7089));
    InMux I__689 (
            .O(N__7102),
            .I(N__7089));
    InMux I__688 (
            .O(N__7101),
            .I(N__7089));
    LocalMux I__687 (
            .O(N__7098),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25));
    LocalMux I__686 (
            .O(N__7089),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25));
    InMux I__685 (
            .O(N__7084),
            .I(N__7081));
    LocalMux I__684 (
            .O(N__7081),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__683 (
            .O(N__7078),
            .I(N__7074));
    InMux I__682 (
            .O(N__7077),
            .I(N__7071));
    LocalMux I__681 (
            .O(N__7074),
            .I(N__7066));
    LocalMux I__680 (
            .O(N__7071),
            .I(N__7066));
    Odrv4 I__679 (
            .O(N__7066),
            .I(un21_beamy_cry_4_c_RNIGUAZ0Z3));
    CascadeMux I__678 (
            .O(N__7063),
            .I(N__7060));
    InMux I__677 (
            .O(N__7060),
            .I(N__7057));
    LocalMux I__676 (
            .O(N__7057),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__675 (
            .O(N__7054),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    CascadeMux I__674 (
            .O(N__7051),
            .I(N__7048));
    InMux I__673 (
            .O(N__7048),
            .I(N__7045));
    LocalMux I__672 (
            .O(N__7045),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICMZ0Z321));
    InMux I__671 (
            .O(N__7042),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__670 (
            .O(N__7039),
            .I(N__7036));
    LocalMux I__669 (
            .O(N__7036),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPMZ0Z1));
    InMux I__668 (
            .O(N__7033),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__667 (
            .O(N__7030),
            .I(N__7027));
    InMux I__666 (
            .O(N__7027),
            .I(N__7024));
    LocalMux I__665 (
            .O(N__7024),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KHZ0Z2));
    InMux I__664 (
            .O(N__7021),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__663 (
            .O(N__7018),
            .I(N__7015));
    LocalMux I__662 (
            .O(N__7015),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__661 (
            .O(N__7012),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__660 (
            .O(N__7009),
            .I(N__7004));
    CascadeMux I__659 (
            .O(N__7008),
            .I(N__7000));
    InMux I__658 (
            .O(N__7007),
            .I(N__6996));
    InMux I__657 (
            .O(N__7004),
            .I(N__6987));
    InMux I__656 (
            .O(N__7003),
            .I(N__6987));
    InMux I__655 (
            .O(N__7000),
            .I(N__6987));
    InMux I__654 (
            .O(N__6999),
            .I(N__6987));
    LocalMux I__653 (
            .O(N__6996),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92));
    LocalMux I__652 (
            .O(N__6987),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92));
    InMux I__651 (
            .O(N__6982),
            .I(N__6979));
    LocalMux I__650 (
            .O(N__6979),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__649 (
            .O(N__6976),
            .I(N__6973));
    LocalMux I__648 (
            .O(N__6973),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__647 (
            .O(N__6970),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__646 (
            .O(N__6967),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01_cascade_));
    CascadeMux I__645 (
            .O(N__6964),
            .I(N__6961));
    InMux I__644 (
            .O(N__6961),
            .I(N__6958));
    LocalMux I__643 (
            .O(N__6958),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__642 (
            .O(N__6955),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__641 (
            .O(N__6952),
            .I(N__6949));
    LocalMux I__640 (
            .O(N__6949),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOLZ0));
    InMux I__639 (
            .O(N__6946),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    CascadeMux I__638 (
            .O(N__6943),
            .I(N__6939));
    InMux I__637 (
            .O(N__6942),
            .I(N__6930));
    InMux I__636 (
            .O(N__6939),
            .I(N__6930));
    InMux I__635 (
            .O(N__6938),
            .I(N__6930));
    InMux I__634 (
            .O(N__6937),
            .I(N__6927));
    LocalMux I__633 (
            .O(N__6930),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01));
    LocalMux I__632 (
            .O(N__6927),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01));
    CascadeMux I__631 (
            .O(N__6922),
            .I(N__6919));
    InMux I__630 (
            .O(N__6919),
            .I(N__6916));
    LocalMux I__629 (
            .O(N__6916),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IGZ0Z1));
    InMux I__628 (
            .O(N__6913),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__627 (
            .O(N__6910),
            .I(N__6907));
    LocalMux I__626 (
            .O(N__6907),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7));
    CascadeMux I__625 (
            .O(N__6904),
            .I(N__6901));
    InMux I__624 (
            .O(N__6901),
            .I(N__6898));
    LocalMux I__623 (
            .O(N__6898),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMGZ0Z1));
    InMux I__622 (
            .O(N__6895),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__621 (
            .O(N__6892),
            .I(N__6889));
    LocalMux I__620 (
            .O(N__6889),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__619 (
            .O(N__6886),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__618 (
            .O(N__6883),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    InMux I__617 (
            .O(N__6880),
            .I(N__6877));
    LocalMux I__616 (
            .O(N__6877),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOGZ0Z53));
    InMux I__615 (
            .O(N__6874),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__614 (
            .O(N__6871),
            .I(N__6868));
    LocalMux I__613 (
            .O(N__6868),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOSZ0));
    InMux I__612 (
            .O(N__6865),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3));
    CascadeMux I__611 (
            .O(N__6862),
            .I(N__6859));
    InMux I__610 (
            .O(N__6859),
            .I(N__6856));
    LocalMux I__609 (
            .O(N__6856),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRSZ0));
    InMux I__608 (
            .O(N__6853),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__607 (
            .O(N__6850),
            .I(N__6847));
    InMux I__606 (
            .O(N__6847),
            .I(N__6844));
    LocalMux I__605 (
            .O(N__6844),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LKZ0));
    InMux I__604 (
            .O(N__6841),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__603 (
            .O(N__6838),
            .I(N__6835));
    LocalMux I__602 (
            .O(N__6835),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_axb_7));
    InMux I__601 (
            .O(N__6832),
            .I(un21_beamy_cry_5));
    InMux I__600 (
            .O(N__6829),
            .I(un21_beamy_cry_6));
    InMux I__599 (
            .O(N__6826),
            .I(un21_beamy_cry_7));
    InMux I__598 (
            .O(N__6823),
            .I(bfn_1_7_0_));
    InMux I__597 (
            .O(N__6820),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__596 (
            .O(N__6817),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__595 (
            .O(N__6814),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__594 (
            .O(N__6811),
            .I(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__593 (
            .O(N__6808),
            .I(un21_beamy_cry_1));
    InMux I__592 (
            .O(N__6805),
            .I(un21_beamy_cry_2));
    InMux I__591 (
            .O(N__6802),
            .I(un21_beamy_cry_3));
    InMux I__590 (
            .O(N__6799),
            .I(un21_beamy_cry_4));
    IoInMux I__589 (
            .O(N__6796),
            .I(N__6793));
    LocalMux I__588 (
            .O(N__6793),
            .I(N__6790));
    Span4Mux_s1_h I__587 (
            .O(N__6790),
            .I(N__6787));
    Span4Mux_h I__586 (
            .O(N__6787),
            .I(N__6784));
    Sp12to4 I__585 (
            .O(N__6784),
            .I(N__6781));
    Odrv12 I__584 (
            .O(N__6781),
            .I(\Clock50MHz.PixelClock ));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(un5_visiblex_cry_7),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(un21_beamy_cry_8),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__6796),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam beamY_5_LC_1_4_0.C_ON=1'b0;
    defparam beamY_5_LC_1_4_0.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_1_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_5_LC_1_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7077),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11877),
            .ce(N__11058),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un5_beamx_4_LC_1_5_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un5_beamx_4_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un5_beamx_4_LC_1_5_0.LUT_INIT=16'b0000000000110011;
    LogicCell40 un114_pixel_1_0_3__un5_beamx_4_LC_1_5_0 (
            .in0(_gnd_net_),
            .in1(N__7590),
            .in2(_gnd_net_),
            .in3(N__7663),
            .lcout(un1_beamy_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_5_LC_1_5_1.C_ON=1'b0;
    defparam beamY_RNI6125_5_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_5_LC_1_5_1.LUT_INIT=16'b1001010101010101;
    LogicCell40 beamY_RNI6125_5_LC_1_5_1 (
            .in0(N__7664),
            .in1(N__12177),
            .in2(N__10632),
            .in3(N__8607),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_4_LC_1_5_7.C_ON=1'b0;
    defparam beamY_RNIBFP3_4_LC_1_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_4_LC_1_5_7.LUT_INIT=16'b0111011110001000;
    LogicCell40 beamY_RNIBFP3_4_LC_1_5_7 (
            .in0(N__10595),
            .in1(N__12178),
            .in2(_gnd_net_),
            .in3(N__8608),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_LC_1_6_0.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_LC_1_6_0.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_LC_1_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_LC_1_6_0 (
            .in0(_gnd_net_),
            .in1(N__14760),
            .in2(N__15008),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(un21_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_RNIAL73_LC_1_6_1.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_1_6_1.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_RNIAL73_LC_1_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_1_c_RNIAL73_LC_1_6_1 (
            .in0(_gnd_net_),
            .in1(N__12208),
            .in2(_gnd_net_),
            .in3(N__6808),
            .lcout(un21_beamy_cry_1_c_RNIALZ0Z73),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_2_c_RNICO83_LC_1_6_2.C_ON=1'b1;
    defparam un21_beamy_cry_2_c_RNICO83_LC_1_6_2.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_2_c_RNICO83_LC_1_6_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_2_c_RNICO83_LC_1_6_2 (
            .in0(_gnd_net_),
            .in1(N__10631),
            .in2(_gnd_net_),
            .in3(N__6805),
            .lcout(un21_beamy_cry_2_c_RNICOZ0Z83),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_4_LC_1_6_3.C_ON=1'b1;
    defparam beamY_4_LC_1_6_3.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_1_6_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_4_LC_1_6_3 (
            .in0(N__10978),
            .in1(N__8620),
            .in2(_gnd_net_),
            .in3(N__6802),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(N__11873),
            .ce(N__11065),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_1_6_4.C_ON=1'b1;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_1_6_4.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_4_c_RNIGUA3_LC_1_6_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_4_c_RNIGUA3_LC_1_6_4 (
            .in0(_gnd_net_),
            .in1(N__7681),
            .in2(_gnd_net_),
            .in3(N__6799),
            .lcout(un21_beamy_cry_4_c_RNIGUAZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_6_LC_1_6_5.C_ON=1'b1;
    defparam beamY_6_LC_1_6_5.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_1_6_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_6_LC_1_6_5 (
            .in0(_gnd_net_),
            .in1(N__7600),
            .in2(_gnd_net_),
            .in3(N__6832),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(N__11873),
            .ce(N__11065),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_1_6_6.C_ON=1'b1;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_1_6_6.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_6_c_RNIK4D3_LC_1_6_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un21_beamy_cry_6_c_RNIK4D3_LC_1_6_6 (
            .in0(_gnd_net_),
            .in1(N__7809),
            .in2(_gnd_net_),
            .in3(N__6829),
            .lcout(un21_beamy_cry_6_c_RNIK4DZ0Z3),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_8_LC_1_6_7.C_ON=1'b1;
    defparam beamY_8_LC_1_6_7.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_1_6_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_1_6_7 (
            .in0(_gnd_net_),
            .in1(N__7922),
            .in2(_gnd_net_),
            .in3(N__6826),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(N__11873),
            .ce(N__11065),
            .sr(_gnd_net_));
    defparam beamY_9_LC_1_7_0.C_ON=1'b0;
    defparam beamY_9_LC_1_7_0.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_1_7_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_9_LC_1_7_0 (
            .in0(N__10954),
            .in1(N__7852),
            .in2(_gnd_net_),
            .in3(N__6823),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11872),
            .ce(N__11068),
            .sr(_gnd_net_));
    defparam beamY_7_LC_1_7_5.C_ON=1'b0;
    defparam beamY_7_LC_1_7_5.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_1_7_5.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_7_LC_1_7_5 (
            .in0(_gnd_net_),
            .in1(N__7203),
            .in2(_gnd_net_),
            .in3(N__10955),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11872),
            .ce(N__11068),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_8_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12804),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOS_LC_1_8_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOS_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOS_LC_1_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOS_LC_1_8_1 (
            .in0(_gnd_net_),
            .in1(N__7306),
            .in2(N__16402),
            .in3(N__6820),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOSZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRS_LC_1_8_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRS_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRS_LC_1_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRS_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(N__7228),
            .in2(N__16407),
            .in3(N__6817),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRSZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LK_LC_1_8_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LK_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LK_LC_1_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LK_LC_1_8_3 (
            .in0(_gnd_net_),
            .in1(N__7213),
            .in2(N__16403),
            .in3(N__6814),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LKZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI8C3M_LC_1_8_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI8C3M_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI8C3M_LC_1_8_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI8C3M_LC_1_8_4 (
            .in0(N__7288),
            .in1(N__6880),
            .in2(N__7336),
            .in3(N__6811),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_1_8_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_1_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_1_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6883),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_1_8_6.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_1_8_6.LUT_INIT=16'b0101010110101010;
    LogicCell40 beamY_RNIHUG2_3_LC_1_8_6 (
            .in0(N__10633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12245),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOG53_LC_1_8_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOG53_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOG53_LC_1_8_7.LUT_INIT=16'b0110011001100110;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOG53_LC_1_8_7 (
            .in0(N__7331),
            .in1(N__7332),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOGZ0Z53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_1_LC_1_9_0.C_ON=1'b1;
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_1_LC_1_9_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_1_LC_1_9_0.LUT_INIT=16'b0000111111110000;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_1_LC_1_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9462),
            .in3(N__10891),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_c5_0_nsZ0Z_1),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOL_LC_1_9_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOL_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOL_LC_1_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOL_LC_1_9_1 (
            .in0(_gnd_net_),
            .in1(N__7289),
            .in2(N__6964),
            .in3(N__6874),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOLZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IG1_LC_1_9_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IG1_LC_1_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IG1_LC_1_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IG1_LC_1_9_2 (
            .in0(_gnd_net_),
            .in1(N__6871),
            .in2(N__7294),
            .in3(N__6865),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IGZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMG1_LC_1_9_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMG1_LC_1_9_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMG1_LC_1_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMG1_LC_1_9_3 (
            .in0(_gnd_net_),
            .in1(N__7293),
            .in2(N__6862),
            .in3(N__6853),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMGZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI70192_LC_1_9_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI70192_LC_1_9_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI70192_LC_1_9_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI70192_LC_1_9_4 (
            .in0(N__6937),
            .in1(N__7267),
            .in2(N__6850),
            .in3(N__6841),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_LC_1_9_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_LC_1_9_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_LC_1_9_5 (
            .in0(N__6838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6970),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01),
            .ltout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_0_LC_1_9_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_0_LC_1_9_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_0_LC_1_9_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_0_LC_1_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6967),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_9_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_9_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12805),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_10_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_10_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_10_0 (
            .in0(_gnd_net_),
            .in1(N__9535),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICM321_LC_1_10_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICM321_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICM321_LC_1_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICM321_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(N__6938),
            .in2(N__7063),
            .in3(N__6955),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICMZ0Z321),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPM1_LC_1_10_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPM1_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPM1_LC_1_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPM1_LC_1_10_2 (
            .in0(_gnd_net_),
            .in1(N__6952),
            .in2(N__6943),
            .in3(N__6946),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPMZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KH2_LC_1_10_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KH2_LC_1_10_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KH2_LC_1_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KH2_LC_1_10_3 (
            .in0(_gnd_net_),
            .in1(N__6942),
            .in2(N__6922),
            .in3(N__6913),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KHZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI1RER4_LC_1_10_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI1RER4_LC_1_10_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI1RER4_LC_1_10_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI1RER4_LC_1_10_4 (
            .in0(N__7007),
            .in1(N__6910),
            .in2(N__6904),
            .in3(N__6895),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_LC_1_10_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_LC_1_10_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_LC_1_10_5 (
            .in0(_gnd_net_),
            .in1(N__6892),
            .in2(_gnd_net_),
            .in3(N__6886),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_10_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_10_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9463),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHGR8_5_LC_1_11_0.C_ON=1'b1;
    defparam beamY_RNIHGR8_5_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIHGR8_5_LC_1_11_0.LUT_INIT=16'b0110011001100110;
    LogicCell40 beamY_RNIHGR8_5_LC_1_11_0 (
            .in0(N__9537),
            .in1(N__9698),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(g0_2_0),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CR2_LC_1_11_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CR2_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CR2_LC_1_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CR2_LC_1_11_1 (
            .in0(_gnd_net_),
            .in1(N__6976),
            .in2(N__7008),
            .in3(N__7054),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CRZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGI3_LC_1_11_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGI3_LC_1_11_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGI3_LC_1_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGI3_LC_1_11_2 (
            .in0(_gnd_net_),
            .in1(N__7003),
            .in2(N__7051),
            .in3(N__7042),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGIZ0Z3),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJ6874_LC_1_11_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJ6874_LC_1_11_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJ6874_LC_1_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJ6874_LC_1_11_3 (
            .in0(_gnd_net_),
            .in1(N__7039),
            .in2(N__7009),
            .in3(N__7033),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJZ0Z6874),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI0RD4A_LC_1_11_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI0RD4A_LC_1_11_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI0RD4A_LC_1_11_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI0RD4A_LC_1_11_4 (
            .in0(N__7107),
            .in1(N__6982),
            .in2(N__7030),
            .in3(N__7021),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_LC_1_11_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_LC_1_11_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_LC_1_11_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_LC_1_11_5 (
            .in0(_gnd_net_),
            .in1(N__7018),
            .in2(_gnd_net_),
            .in3(N__7012),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_0_LC_1_11_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_0_LC_1_11_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_0_LC_1_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_0_LC_1_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6999),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_11_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_11_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9536),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_12_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_12_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_12_0 (
            .in0(_gnd_net_),
            .in1(N__8522),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_12_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEG5_LC_1_12_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEG5_LC_1_12_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEG5_LC_1_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEG5_LC_1_12_1 (
            .in0(_gnd_net_),
            .in1(N__7102),
            .in2(N__7117),
            .in3(N__7162),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEGZ0Z5),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87V68_LC_1_12_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87V68_LC_1_12_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87V68_LC_1_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87V68_LC_1_12_2 (
            .in0(_gnd_net_),
            .in1(N__7159),
            .in2(N__7108),
            .in3(N__7153),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87VZ0Z68),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05U8_LC_1_12_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05U8_LC_1_12_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05U8_LC_1_12_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05U8_LC_1_12_3 (
            .in0(_gnd_net_),
            .in1(N__7106),
            .in2(N__7150),
            .in3(N__7141),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05UZ0Z8),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIE5N0K_LC_1_12_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIE5N0K_LC_1_12_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIE5N0K_LC_1_12_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIE5N0K_LC_1_12_4 (
            .in0(N__7386),
            .in1(N__7084),
            .in2(N__7138),
            .in3(N__7129),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDA_LC_1_12_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDA_LC_1_12_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDA_LC_1_12_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDA_LC_1_12_5 (
            .in0(_gnd_net_),
            .in1(N__7126),
            .in2(_gnd_net_),
            .in3(N__7120),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_12_6.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_12_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9699),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_0_LC_1_12_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_0_LC_1_12_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_0_LC_1_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_0_LC_1_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7101),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_5_LC_2_4_0.C_ON=1'b0;
    defparam beamY_fast_5_LC_2_4_0.SEQ_MODE=4'b1000;
    defparam beamY_fast_5_LC_2_4_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_5_LC_2_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7078),
            .lcout(beamY_fastZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11880),
            .ce(N__11057),
            .sr(_gnd_net_));
    defparam beamY_2_LC_2_5_1.C_ON=1'b0;
    defparam beamY_2_LC_2_5_1.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_2_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_2_LC_2_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7174),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11878),
            .ce(N__11067),
            .sr(_gnd_net_));
    defparam beamY_3_LC_2_5_3.C_ON=1'b0;
    defparam beamY_3_LC_2_5_3.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_2_5_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 beamY_3_LC_2_5_3 (
            .in0(_gnd_net_),
            .in1(N__10974),
            .in2(_gnd_net_),
            .in3(N__7243),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11878),
            .ce(N__11067),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIVDP7_7_LC_2_5_5.C_ON=1'b0;
    defparam beamY_fast_RNIVDP7_7_LC_2_5_5.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIVDP7_7_LC_2_5_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 beamY_fast_RNIVDP7_7_LC_2_5_5 (
            .in0(N__7911),
            .in1(N__7588),
            .in2(N__7192),
            .in3(N__7662),
            .lcout(un5_visibley_ac0_11_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_7_LC_2_5_6.C_ON=1'b0;
    defparam beamY_fast_7_LC_2_5_6.SEQ_MODE=4'b1000;
    defparam beamY_fast_7_LC_2_5_6.LUT_INIT=16'b0100010001000100;
    LogicCell40 beamY_fast_7_LC_2_5_6 (
            .in0(N__10975),
            .in1(N__7204),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11878),
            .ce(N__11067),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIEP79_5_LC_2_5_7.C_ON=1'b0;
    defparam beamY_fast_RNIEP79_5_LC_2_5_7.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIEP79_5_LC_2_5_7.LUT_INIT=16'b1111111111101110;
    LogicCell40 beamY_fast_RNIEP79_5_LC_2_5_7 (
            .in0(N__7191),
            .in1(N__7180),
            .in2(_gnd_net_),
            .in3(N__7589),
            .lcout(un5_visibley_c6_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIP81D_7_LC_2_6_0.C_ON=1'b0;
    defparam beamY_RNIP81D_7_LC_2_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIP81D_7_LC_2_6_0.LUT_INIT=16'b1000011111110000;
    LogicCell40 beamY_RNIP81D_7_LC_2_6_0 (
            .in0(N__8601),
            .in1(N__7994),
            .in2(N__7810),
            .in3(N__7955),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_2_LC_2_6_2.C_ON=1'b0;
    defparam beamY_fast_2_LC_2_6_2.SEQ_MODE=4'b1000;
    defparam beamY_fast_2_LC_2_6_2.LUT_INIT=16'b1100110011001100;
    LogicCell40 beamY_fast_2_LC_2_6_2 (
            .in0(_gnd_net_),
            .in1(N__7173),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11875),
            .ce(N__11066),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI35GA_0_2_LC_2_6_3.C_ON=1'b0;
    defparam beamY_fast_RNI35GA_0_2_LC_2_6_3.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI35GA_0_2_LC_2_6_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 beamY_fast_RNI35GA_0_2_LC_2_6_3 (
            .in0(N__7708),
            .in1(N__7906),
            .in2(N__7638),
            .in3(N__8599),
            .lcout(un5_visibley_ac0_11_d),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNI35GA_2_LC_2_6_4.C_ON=1'b0;
    defparam beamY_fast_RNI35GA_2_LC_2_6_4.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNI35GA_2_LC_2_6_4.LUT_INIT=16'b1000011100001111;
    LogicCell40 beamY_fast_RNI35GA_2_LC_2_6_4 (
            .in0(N__8600),
            .in1(N__7633),
            .in2(N__7923),
            .in3(N__7709),
            .lcout(),
            .ltout(beamY_fast_RNI35GAZ0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFJ0L_8_LC_2_6_5.C_ON=1'b0;
    defparam beamY_RNIFJ0L_8_LC_2_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIFJ0L_8_LC_2_6_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 beamY_RNIFJ0L_8_LC_2_6_5 (
            .in0(N__7252),
            .in1(_gnd_net_),
            .in2(N__7246),
            .in3(N__7910),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_3_LC_2_6_6.C_ON=1'b0;
    defparam beamY_fast_3_LC_2_6_6.SEQ_MODE=4'b1000;
    defparam beamY_fast_3_LC_2_6_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_fast_3_LC_2_6_6 (
            .in0(_gnd_net_),
            .in1(N__7242),
            .in2(_gnd_net_),
            .in3(N__10976),
            .lcout(beamY_fastZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11875),
            .ce(N__11066),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_7_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_7_0 (
            .in0(_gnd_net_),
            .in1(N__12538),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_2_7_1.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_2_7_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_2_7_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_2_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7231),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI19IJ_9_LC_2_7_3.C_ON=1'b0;
    defparam beamY_RNI19IJ_9_LC_2_7_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI19IJ_9_LC_2_7_3.LUT_INIT=16'b1010101010011001;
    LogicCell40 beamY_RNI19IJ_9_LC_2_7_3 (
            .in0(N__7844),
            .in1(N__7758),
            .in2(_gnd_net_),
            .in3(N__7743),
            .lcout(chary_if_generate_plus_mult1_un33_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un8_beamylto4_0_LC_2_7_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un8_beamylto4_0_LC_2_7_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un8_beamylto4_0_LC_2_7_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 un114_pixel_1_0_3__un8_beamylto4_0_LC_2_7_5 (
            .in0(N__7710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7634),
            .lcout(un5_visibley_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_8_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_8_0 (
            .in0(_gnd_net_),
            .in1(N__12654),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2L_LC_2_8_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2L_LC_2_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2L_LC_2_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2L_LC_2_8_1 (
            .in0(_gnd_net_),
            .in1(N__7300),
            .in2(N__16383),
            .in3(N__7222),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2LZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RC_LC_2_8_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RC_LC_2_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RC_LC_2_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RC_LC_2_8_2 (
            .in0(_gnd_net_),
            .in1(N__7219),
            .in2(N__16384),
            .in3(N__7207),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RCZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOI1_LC_2_8_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOI1_LC_2_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOI1_LC_2_8_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOI1_LC_2_8_3 (
            .in0(_gnd_net_),
            .in1(N__16355),
            .in2(_gnd_net_),
            .in3(N__7318),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_LC_2_8_4.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_LC_2_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_LC_2_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_LC_2_8_4 (
            .in0(_gnd_net_),
            .in1(N__7315),
            .in2(_gnd_net_),
            .in3(N__7309),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFJ0L_0_8_LC_2_8_5.C_ON=1'b0;
    defparam beamY_RNIFJ0L_0_8_LC_2_8_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIFJ0L_0_8_LC_2_8_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 beamY_RNIFJ0L_0_8_LC_2_8_5 (
            .in0(N__12655),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_RNIFJ0L_0Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI19IJ_0_9_LC_2_8_7.C_ON=1'b0;
    defparam beamY_RNI19IJ_0_9_LC_2_8_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI19IJ_0_9_LC_2_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 beamY_RNI19IJ_0_9_LC_2_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12539),
            .lcout(beamY_RNI19IJ_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_0_LC_2_9_1.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_0_LC_2_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_0_LC_2_9_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_0_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7287),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_9_2.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_9_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_9_2 (
            .in0(N__7484),
            .in1(N__16401),
            .in2(_gnd_net_),
            .in3(N__12246),
            .lcout(beamY_i_2),
            .ltout(beamY_i_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_1_LC_2_9_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_1_LC_2_9_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_1_LC_2_9_3.LUT_INIT=16'b0001100010001000;
    LogicCell40 un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_1_LC_2_9_3 (
            .in0(N__7461),
            .in1(N__7437),
            .in2(N__7261),
            .in3(N__7346),
            .lcout(),
            .ltout(un114_pixel_1_0_3__chessboardpixel_un200_pixellto4Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_LC_2_9_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_LC_2_9_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_LC_2_9_4.LUT_INIT=16'b1000000001000000;
    LogicCell40 un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_LC_2_9_4 (
            .in0(N__7347),
            .in1(N__15013),
            .in2(N__7258),
            .in3(N__7485),
            .lcout(),
            .ltout(chessboardpixel_un200_pixellt10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto10_1_LC_2_9_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto10_1_LC_2_9_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__chessboardpixel_un200_pixellto10_1_LC_2_9_5.LUT_INIT=16'b0000011000000101;
    LogicCell40 un114_pixel_1_0_3__chessboardpixel_un200_pixellto10_1_LC_2_9_5 (
            .in0(N__7417),
            .in1(N__7492),
            .in2(N__7255),
            .in3(N__7348),
            .lcout(),
            .ltout(chessboardpixel_un200_pixel_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__Pixel_3_sqmuxa_0_LC_2_9_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__Pixel_3_sqmuxa_0_LC_2_9_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__Pixel_3_sqmuxa_0_LC_2_9_6.LUT_INIT=16'b0000110011000000;
    LogicCell40 un114_pixel_1_0_3__Pixel_3_sqmuxa_0_LC_2_9_6 (
            .in0(_gnd_net_),
            .in1(N__12118),
            .in2(N__7495),
            .in3(N__7558),
            .lcout(un114_pixel_1_0_3__Pixel_3_sqmuxaZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIMR0FR_LC_2_9_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIMR0FR_LC_2_9_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIMR0FR_LC_2_9_7.LUT_INIT=16'b1111111110111011;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIMR0FR_LC_2_9_7 (
            .in0(N__7462),
            .in1(N__7483),
            .in2(_gnd_net_),
            .in3(N__7438),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_10_0.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_10_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7486),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81B_LC_2_10_1.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81B_LC_2_10_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81B_LC_2_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81B_LC_2_10_1 (
            .in0(_gnd_net_),
            .in1(N__7552),
            .in2(N__7395),
            .in3(N__7453),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81BZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODG_LC_2_10_2.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODG_LC_2_10_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODG_LC_2_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODG_LC_2_10_2 (
            .in0(_gnd_net_),
            .in1(N__7391),
            .in2(N__7450),
            .in3(N__7429),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODGZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4J_LC_2_10_3.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4J_LC_2_10_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4J_LC_2_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4J_LC_2_10_3 (
            .in0(_gnd_net_),
            .in1(N__7426),
            .in2(N__7396),
            .in3(N__7411),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4JZ0),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_10_4.C_ON=1'b1;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_10_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_10_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(N__7366),
            .in2(N__7408),
            .in3(N__7387),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGK_LC_2_10_5.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGK_LC_2_10_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGK_LC_2_10_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGK_LC_2_10_5 (
            .in0(_gnd_net_),
            .in1(N__7360),
            .in2(_gnd_net_),
            .in3(N__7351),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGKZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_LC_2_10_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_LC_2_10_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_LC_2_10_6.LUT_INIT=16'b1000001010010010;
    LogicCell40 un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_LC_2_10_6 (
            .in0(N__7501),
            .in1(N__7513),
            .in2(N__7528),
            .in3(N__11544),
            .lcout(chessboardpixel_un174_pixel_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_10_7.C_ON=1'b0;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_10_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8523),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_2_11_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_2_11_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_2_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_2_11_0 (
            .in0(_gnd_net_),
            .in1(N__11547),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJ5_LC_2_11_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJ5_LC_2_11_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJ5_LC_2_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJ5_LC_2_11_1 (
            .in0(_gnd_net_),
            .in1(N__7539),
            .in2(N__9043),
            .in3(N__7546),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJZ0Z5),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAEC_LC_2_11_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAEC_LC_2_11_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAEC_LC_2_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAEC_LC_2_11_2 (
            .in0(_gnd_net_),
            .in1(N__8203),
            .in2(N__8248),
            .in3(N__7543),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_2_11_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_2_11_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_2_11_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_2_11_3 (
            .in0(N__8202),
            .in1(N__7540),
            .in2(N__8233),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHF_LC_2_11_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHF_LC_2_11_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHF_LC_2_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHF_LC_2_11_4 (
            .in0(_gnd_net_),
            .in1(N__8218),
            .in2(_gnd_net_),
            .in3(N__7531),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHFZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_1_LC_2_11_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_1_LC_2_11_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_1_LC_2_11_6.LUT_INIT=16'b0101011100010101;
    LogicCell40 un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_1_LC_2_11_6 (
            .in0(N__7519),
            .in1(N__7512),
            .in2(N__13612),
            .in3(N__11548),
            .lcout(un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKHPCA1_4_LC_4_3_5.C_ON=1'b0;
    defparam beamY_RNIKHPCA1_4_LC_4_3_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIKHPCA1_4_LC_4_3_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNIKHPCA1_4_LC_4_3_5 (
            .in0(N__9765),
            .in1(N__9298),
            .in2(_gnd_net_),
            .in3(N__9933),
            .lcout(beamY_RNIKHPCA1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISKOB_5_LC_4_5_0.C_ON=1'b0;
    defparam beamY_RNISKOB_5_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNISKOB_5_LC_4_5_0.LUT_INIT=16'b1010101010010101;
    LogicCell40 beamY_RNISKOB_5_LC_4_5_0 (
            .in0(N__7608),
            .in1(N__8641),
            .in2(N__8008),
            .in3(N__7682),
            .lcout(chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un1_beamylto9_0_LC_4_5_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un1_beamylto9_0_LC_4_5_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un1_beamylto9_0_LC_4_5_3.LUT_INIT=16'b0000000000110011;
    LogicCell40 un114_pixel_1_0_3__un1_beamylto9_0_LC_4_5_3 (
            .in0(_gnd_net_),
            .in1(N__10641),
            .in2(_gnd_net_),
            .in3(N__7825),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un1_beamylto9Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un1_beamylto9_3_0_LC_4_5_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un1_beamylto9_3_0_LC_4_5_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un1_beamylto9_3_0_LC_4_5_4.LUT_INIT=16'b0000000001110000;
    LogicCell40 un114_pixel_1_0_3__un1_beamylto9_3_0_LC_4_5_4 (
            .in0(N__14994),
            .in1(N__12216),
            .in2(N__7768),
            .in3(N__8642),
            .lcout(un114_pixel_1_0_3__un1_beamylto9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_1_3_LC_4_5_6.C_ON=1'b0;
    defparam beamY_RNIHUG2_1_3_LC_4_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_1_3_LC_4_5_6.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIHUG2_1_3_LC_4_5_6 (
            .in0(N__10640),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12215),
            .lcout(un4_beamylt6),
            .ltout(un4_beamylt6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_beamylto6_LC_4_5_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_beamylto6_LC_4_5_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_beamylto6_LC_4_5_7.LUT_INIT=16'b0000100000000000;
    LogicCell40 un114_pixel_1_0_3__un4_beamylto6_LC_4_5_7 (
            .in0(N__7683),
            .in1(N__7609),
            .in2(N__7765),
            .in3(N__8643),
            .lcout(un4_beamylt8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDO3I_9_LC_4_6_0.C_ON=1'b0;
    defparam beamY_RNIDO3I_9_LC_4_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIDO3I_9_LC_4_6_0.LUT_INIT=16'b1011110101010101;
    LogicCell40 beamY_RNIDO3I_9_LC_4_6_0 (
            .in0(N__7871),
            .in1(N__7823),
            .in2(N__8038),
            .in3(N__7924),
            .lcout(beamY_RNIDO3IZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGSI81_9_LC_4_6_2.C_ON=1'b0;
    defparam beamY_RNIGSI81_9_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIGSI81_9_LC_4_6_2.LUT_INIT=16'b0101000001100000;
    LogicCell40 beamY_RNIGSI81_9_LC_4_6_2 (
            .in0(N__7870),
            .in1(N__7762),
            .in2(N__12685),
            .in3(N__7747),
            .lcout(chary_if_generate_plus_mult1_un40_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un1_beamylto9_LC_4_6_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un1_beamylto9_LC_4_6_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un1_beamylto9_LC_4_6_4.LUT_INIT=16'b0000000001000000;
    LogicCell40 un114_pixel_1_0_3__un1_beamylto9_LC_4_6_4 (
            .in0(N__7872),
            .in1(N__7978),
            .in2(N__7726),
            .in3(N__7925),
            .lcout(un1_beamylto9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIM4P7_2_LC_4_6_5.C_ON=1'b0;
    defparam beamY_fast_RNIM4P7_2_LC_4_6_5.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIM4P7_2_LC_4_6_5.LUT_INIT=16'b1111111111101100;
    LogicCell40 beamY_fast_RNIM4P7_2_LC_4_6_5 (
            .in0(N__8629),
            .in1(N__7606),
            .in2(N__7717),
            .in3(N__7689),
            .lcout(),
            .ltout(beamY_fast_RNIM4P7Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIJP9E_3_LC_4_6_6.C_ON=1'b0;
    defparam beamY_fast_RNIJP9E_3_LC_4_6_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIJP9E_3_LC_4_6_6.LUT_INIT=16'b1111001111100010;
    LogicCell40 beamY_fast_RNIJP9E_3_LC_4_6_6 (
            .in0(N__7690),
            .in1(N__7639),
            .in2(N__7612),
            .in3(N__7607),
            .lcout(un5_visibley_c5),
            .ltout(un5_visibley_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0A5O1_7_LC_4_6_7.C_ON=1'b0;
    defparam beamY_RNI0A5O1_7_LC_4_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI0A5O1_7_LC_4_6_7.LUT_INIT=16'b0011001110110111;
    LogicCell40 beamY_RNI0A5O1_7_LC_4_6_7 (
            .in0(N__7824),
            .in1(N__12665),
            .in2(N__8029),
            .in3(N__12581),
            .lcout(chary_if_generate_plus_mult1_un40_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un5_beamx_5_LC_4_7_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un5_beamx_5_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un5_beamx_5_LC_4_7_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_1_0_3__un5_beamx_5_LC_4_7_0 (
            .in0(N__7819),
            .in1(N__15007),
            .in2(N__8659),
            .in3(N__7874),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un5_beamxZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un5_beamx_LC_4_7_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un5_beamx_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un5_beamx_LC_4_7_1.LUT_INIT=16'b0000000010000000;
    LogicCell40 un114_pixel_1_0_3__un5_beamx_LC_4_7_1 (
            .in0(N__8645),
            .in1(N__7977),
            .in2(N__8026),
            .in3(N__7939),
            .lcout(un5_beamx_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_1_0_LC_4_7_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_1_0_LC_4_7_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_1_0_LC_4_7_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 un114_pixel_1_0_3__g0_1_0_LC_4_7_2 (
            .in0(_gnd_net_),
            .in1(N__7875),
            .in2(_gnd_net_),
            .in3(N__7938),
            .lcout(),
            .ltout(un114_pixel_1_0_3__g0_1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_3_LC_4_7_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_3_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_3_LC_4_7_3.LUT_INIT=16'b0000000010000000;
    LogicCell40 un114_pixel_1_0_3__g0_3_LC_4_7_3 (
            .in0(N__7976),
            .in1(N__8563),
            .in2(N__8023),
            .in3(N__7818),
            .lcout(un1_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_beamylto9_LC_4_7_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_beamylto9_LC_4_7_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_beamylto9_LC_4_7_4.LUT_INIT=16'b1100110011001000;
    LogicCell40 un114_pixel_1_0_3__un4_beamylto9_LC_4_7_4 (
            .in0(N__7816),
            .in1(N__7873),
            .in2(N__8020),
            .in3(N__7936),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un8_beamylto9_1_LC_4_7_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un8_beamylto9_1_LC_4_7_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un8_beamylto9_1_LC_4_7_6.LUT_INIT=16'b0100010011001100;
    LogicCell40 un114_pixel_1_0_3__un8_beamylto9_1_LC_4_7_6 (
            .in0(N__8004),
            .in1(N__7975),
            .in2(_gnd_net_),
            .in3(N__8644),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un8_beamylto9Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un8_beamylto9_LC_4_7_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un8_beamylto9_LC_4_7_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un8_beamylto9_LC_4_7_7.LUT_INIT=16'b0000000000010000;
    LogicCell40 un114_pixel_1_0_3__un8_beamylto9_LC_4_7_7 (
            .in0(N__7937),
            .in1(N__7876),
            .in2(N__7828),
            .in3(N__7817),
            .lcout(un8_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_8_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_8_1.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_8_1 (
            .in0(N__9764),
            .in1(N__8064),
            .in2(N__8548),
            .in3(N__8157),
            .lcout(if_generate_plus_mult1_un75_sum_axbxc3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un54_sum_c5_LC_4_8_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un54_sum_c5_LC_4_8_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un54_sum_c5_LC_4_8_2.LUT_INIT=16'b1011001001100100;
    LogicCell40 row_1_if_generate_plus_mult1_un54_sum_c5_LC_4_8_2 (
            .in0(N__12816),
            .in1(N__12687),
            .in2(N__9460),
            .in3(N__12591),
            .lcout(row_1_if_generate_plus_mult1_un54_sum_cZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_4_8_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_4_8_3.LUT_INIT=16'b1110000110000111;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_4_8_3 (
            .in0(N__8080),
            .in1(N__8050),
            .in2(N__12417),
            .in3(N__12437),
            .lcout(row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_LC_4_8_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_LC_4_8_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_c5_LC_4_8_5.LUT_INIT=16'b1110101110000010;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_c5_LC_4_8_5 (
            .in0(N__8079),
            .in1(N__8065),
            .in2(N__8158),
            .in3(N__8049),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_cZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_c4_LC_4_8_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_c4_LC_4_8_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_c4_LC_4_8_6.LUT_INIT=16'b0110000011110110;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_c4_LC_4_8_6 (
            .in0(N__8063),
            .in1(N__8153),
            .in2(N__8547),
            .in3(N__9763),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_cZ0Z4),
            .ltout(row_1_if_generate_plus_mult1_un75_sum_cZ0Z4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_8_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_8_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_8_7.LUT_INIT=16'b0110101010101001;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_8_7 (
            .in0(N__12410),
            .in1(N__8048),
            .in2(N__8071),
            .in3(N__12436),
            .lcout(if_generate_plus_mult1_un75_sum_axbxc5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_LC_4_9_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_LC_4_9_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_c4_LC_4_9_0.LUT_INIT=16'b1010101010111011;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_c4_LC_4_9_0 (
            .in0(N__8131),
            .in1(N__10877),
            .in2(_gnd_net_),
            .in3(N__9445),
            .lcout(),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_9_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_9_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_9_1.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_9_1 (
            .in0(N__10878),
            .in1(N__8125),
            .in2(N__8068),
            .in3(N__12721),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1),
            .ltout(row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_LC_4_9_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_LC_4_9_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc5_LC_4_9_2.LUT_INIT=16'b0000111111110000;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc5_LC_4_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8053),
            .in3(N__8152),
            .lcout(if_generate_plus_mult1_un68_sum_axbxc5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc3_LC_4_9_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc3_LC_4_9_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_axbxc3_LC_4_9_3.LUT_INIT=16'b0110011010011001;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_axbxc3_LC_4_9_3 (
            .in0(N__9762),
            .in1(N__12722),
            .in2(_gnd_net_),
            .in3(N__9591),
            .lcout(if_generate_plus_mult1_un68_sum_axbxc3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc3_LC_4_9_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc3_LC_4_9_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un54_sum_axbxc3_LC_4_9_5.LUT_INIT=16'b0110100111010010;
    LogicCell40 row_1_if_generate_plus_mult1_un54_sum_axbxc3_LC_4_9_5 (
            .in0(N__12812),
            .in1(N__12679),
            .in2(N__9461),
            .in3(N__12592),
            .lcout(if_generate_plus_mult1_un54_sum_axbxc3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_LC_4_9_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_LC_4_9_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_LC_4_9_6.LUT_INIT=16'b0101111001011000;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_LC_4_9_6 (
            .in0(N__9590),
            .in1(N__8095),
            .in2(N__8170),
            .in3(N__9761),
            .lcout(row_1_if_generate_plus_mult1_un68_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_10_0.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_10_0.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_10_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_10_0 (
            .in0(N__9449),
            .in1(N__10883),
            .in2(_gnd_net_),
            .in3(N__9571),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_1_0_LC_4_10_1.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_1_0_LC_4_10_1.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_1_0_LC_4_10_1.LUT_INIT=16'b0100100111011011;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_axbxc5_1_0_LC_4_10_1 (
            .in0(N__12811),
            .in1(N__12689),
            .in2(N__12599),
            .in3(N__9448),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_10_2.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_10_2.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_10_2 (
            .in0(_gnd_net_),
            .in1(N__8110),
            .in2(N__8134),
            .in3(N__10882),
            .lcout(if_generate_plus_mult1_un61_sum_axbxc5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_5_LC_4_10_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_5_LC_4_10_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_5_LC_4_10_3.LUT_INIT=16'b0100010010001000;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_5_LC_4_10_3 (
            .in0(N__10879),
            .in1(N__9570),
            .in2(_gnd_net_),
            .in3(N__9446),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_10_4.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_10_4.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_10_4.LUT_INIT=16'b1111111011101010;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_10_4 (
            .in0(N__8089),
            .in1(N__8124),
            .in2(N__8113),
            .in3(N__10880),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_c5),
            .ltout(row_1_if_generate_plus_mult1_un61_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_bm_LC_4_10_5.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_bm_LC_4_10_5.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un68_sum_c5_0_bm_LC_4_10_5.LUT_INIT=16'b0101101010100101;
    LogicCell40 row_1_if_generate_plus_mult1_un68_sum_c5_0_bm_LC_4_10_5 (
            .in0(N__10881),
            .in1(_gnd_net_),
            .in2(N__8104),
            .in3(N__8101),
            .lcout(if_generate_plus_mult1_un68_sum_c5_0_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_c_0_LC_4_10_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_c_0_LC_4_10_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un61_sum_ac0_7_c_0_LC_4_10_7.LUT_INIT=16'b0000000010010010;
    LogicCell40 row_1_if_generate_plus_mult1_un61_sum_ac0_7_c_0_LC_4_10_7 (
            .in0(N__12810),
            .in1(N__12688),
            .in2(N__12598),
            .in3(N__9447),
            .lcout(row_1_if_generate_plus_mult1_un61_sum_ac0_7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_4_11_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_4_11_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_4_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_4_11_0 (
            .in0(_gnd_net_),
            .in1(N__11656),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KC4_LC_4_11_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KC4_LC_4_11_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KC4_LC_4_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KC4_LC_4_11_1 (
            .in0(_gnd_net_),
            .in1(N__8184),
            .in2(N__9052),
            .in3(N__8236),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KCZ0Z4),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGS6_LC_4_11_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGS6_LC_4_11_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGS6_LC_4_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGS6_LC_4_11_2 (
            .in0(_gnd_net_),
            .in1(N__13957),
            .in2(N__13915),
            .in3(N__8221),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGSZ0Z6),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI88ODF_LC_4_11_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI88ODF_LC_4_11_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI88ODF_LC_4_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI88ODF_LC_4_11_3 (
            .in0(N__8201),
            .in1(N__8185),
            .in2(N__13945),
            .in3(N__8209),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3U7_LC_4_11_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3U7_LC_4_11_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3U7_LC_4_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3U7_LC_4_11_4 (
            .in0(_gnd_net_),
            .in1(N__13930),
            .in2(_gnd_net_),
            .in3(N__8206),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_0_LC_4_11_7.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_0_LC_4_11_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_0_LC_4_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_0_LC_4_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13911),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_cry_1_c_LC_4_13_0.C_ON=1'b1;
    defparam counter_cry_1_c_LC_4_13_0.SEQ_MODE=4'b0000;
    defparam counter_cry_1_c_LC_4_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 counter_cry_1_c_LC_4_13_0 (
            .in0(_gnd_net_),
            .in1(N__8263),
            .in2(N__8350),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(counter_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNO_0_2_LC_4_13_1.C_ON=1'b1;
    defparam counter_RNO_0_2_LC_4_13_1.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_2_LC_4_13_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_2_LC_4_13_1 (
            .in0(_gnd_net_),
            .in1(N__8320),
            .in2(_gnd_net_),
            .in3(N__8176),
            .lcout(counter_30),
            .ltout(),
            .carryin(counter_cry_1),
            .carryout(counter_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNO_0_3_LC_4_13_2.C_ON=1'b1;
    defparam counter_RNO_0_3_LC_4_13_2.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_3_LC_4_13_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_3_LC_4_13_2 (
            .in0(_gnd_net_),
            .in1(N__8366),
            .in2(_gnd_net_),
            .in3(N__8173),
            .lcout(counter_29),
            .ltout(),
            .carryin(counter_cry_2),
            .carryout(counter_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNO_0_4_LC_4_13_3.C_ON=1'b1;
    defparam counter_RNO_0_4_LC_4_13_3.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_4_LC_4_13_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 counter_RNO_0_4_LC_4_13_3 (
            .in0(_gnd_net_),
            .in1(N__8937),
            .in2(_gnd_net_),
            .in3(N__8293),
            .lcout(counter_28),
            .ltout(),
            .carryin(counter_cry_3),
            .carryout(counter_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNO_0_5_LC_4_13_4.C_ON=1'b0;
    defparam counter_RNO_0_5_LC_4_13_4.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_5_LC_4_13_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 counter_RNO_0_5_LC_4_13_4 (
            .in0(_gnd_net_),
            .in1(N__9021),
            .in2(_gnd_net_),
            .in3(N__8290),
            .lcout(counter_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNI6R5D_0_LC_4_13_5.C_ON=1'b0;
    defparam counter_RNI6R5D_0_LC_4_13_5.SEQ_MODE=4'b0000;
    defparam counter_RNI6R5D_0_LC_4_13_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 counter_RNI6R5D_0_LC_4_13_5 (
            .in0(N__8264),
            .in1(N__8368),
            .in2(N__8349),
            .in3(N__8319),
            .lcout(slaveselect_1_0_4),
            .ltout(slaveselect_1_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIVUOJ_5_LC_4_13_6.C_ON=1'b0;
    defparam counter_RNIVUOJ_5_LC_4_13_6.SEQ_MODE=4'b0000;
    defparam counter_RNIVUOJ_5_LC_4_13_6.LUT_INIT=16'b0000000011110101;
    LogicCell40 counter_RNIVUOJ_5_LC_4_13_6 (
            .in0(N__8938),
            .in1(_gnd_net_),
            .in2(N__8287),
            .in3(N__9022),
            .lcout(un3_slaveselect),
            .ltout(un3_slaveselect_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_2_LC_4_13_7.C_ON=1'b0;
    defparam counter_2_LC_4_13_7.SEQ_MODE=4'b1000;
    defparam counter_2_LC_4_13_7.LUT_INIT=16'b1000000011000100;
    LogicCell40 counter_2_LC_4_13_7 (
            .in0(N__8900),
            .in1(N__8284),
            .in2(N__8278),
            .in3(N__8858),
            .lcout(counterZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14325),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_3_LC_4_14_1.C_ON=1'b0;
    defparam counter_3_LC_4_14_1.SEQ_MODE=4'b1000;
    defparam counter_3_LC_4_14_1.LUT_INIT=16'b1100010100000000;
    LogicCell40 counter_3_LC_4_14_1 (
            .in0(N__8851),
            .in1(N__8971),
            .in2(N__8911),
            .in3(N__8275),
            .lcout(counterZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14326),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNO_0_1_LC_4_14_3.C_ON=1'b0;
    defparam counter_RNO_0_1_LC_4_14_3.SEQ_MODE=4'b0000;
    defparam counter_RNO_0_1_LC_4_14_3.LUT_INIT=16'b1010010101011010;
    LogicCell40 counter_RNO_0_1_LC_4_14_3 (
            .in0(N__8348),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8265),
            .lcout(),
            .ltout(counter_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_1_LC_4_14_4.C_ON=1'b0;
    defparam counter_1_LC_4_14_4.SEQ_MODE=4'b1000;
    defparam counter_1_LC_4_14_4.LUT_INIT=16'b1000000010110000;
    LogicCell40 counter_1_LC_4_14_4 (
            .in0(N__8970),
            .in1(N__8907),
            .in2(N__8269),
            .in3(N__8852),
            .lcout(counterZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14326),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_0_LC_4_14_5.C_ON=1'b0;
    defparam counter_0_LC_4_14_5.SEQ_MODE=4'b1000;
    defparam counter_0_LC_4_14_5.LUT_INIT=16'b0000000011000101;
    LogicCell40 counter_0_LC_4_14_5 (
            .in0(N__8850),
            .in1(N__8969),
            .in2(N__8910),
            .in3(N__8266),
            .lcout(counterZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14326),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIKUI6_1_LC_4_14_6.C_ON=1'b0;
    defparam counter_RNIKUI6_1_LC_4_14_6.SEQ_MODE=4'b0000;
    defparam counter_RNIKUI6_1_LC_4_14_6.LUT_INIT=16'b0000000000110011;
    LogicCell40 counter_RNIKUI6_1_LC_4_14_6 (
            .in0(_gnd_net_),
            .in1(N__8367),
            .in2(_gnd_net_),
            .in3(N__8347),
            .lcout(),
            .ltout(un1_counterlto3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNINHFG_2_LC_4_14_7.C_ON=1'b0;
    defparam counter_RNINHFG_2_LC_4_14_7.SEQ_MODE=4'b0000;
    defparam counter_RNINHFG_2_LC_4_14_7.LUT_INIT=16'b1000100000001000;
    LogicCell40 counter_RNINHFG_2_LC_4_14_7 (
            .in0(N__8939),
            .in1(N__9023),
            .in2(N__8323),
            .in3(N__8318),
            .lcout(un1_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_2_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_2_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_2_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIS857F2_4_LC_5_3_0.C_ON=1'b0;
    defparam beamY_RNIS857F2_4_LC_5_3_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIS857F2_4_LC_5_3_0.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIS857F2_4_LC_5_3_0 (
            .in0(N__9934),
            .in1(N__10045),
            .in2(N__9783),
            .in3(N__9296),
            .lcout(),
            .ltout(g0_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJU3OQ8_4_LC_5_3_1.C_ON=1'b0;
    defparam beamY_RNIJU3OQ8_4_LC_5_3_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIJU3OQ8_4_LC_5_3_1.LUT_INIT=16'b0101101001101001;
    LogicCell40 beamY_RNIJU3OQ8_4_LC_5_3_1 (
            .in0(N__9361),
            .in1(N__9859),
            .in2(N__8302),
            .in3(N__9257),
            .lcout(g0_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUAPPF4_0_3_LC_5_4_0.C_ON=1'b0;
    defparam beamY_RNIUAPPF4_0_3_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIUAPPF4_0_3_LC_5_4_0.LUT_INIT=16'b0100110110001110;
    LogicCell40 beamY_RNIUAPPF4_0_3_LC_5_4_0 (
            .in0(N__10048),
            .in1(N__8546),
            .in2(N__9782),
            .in3(N__8299),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_1_LC_5_4_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_1_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_1_LC_5_4_1.LUT_INIT=16'b0111111010000001;
    LogicCell40 un114_pixel_1_0_3__g0_1_LC_5_4_1 (
            .in0(N__8434),
            .in1(N__9081),
            .in2(N__8377),
            .in3(N__9358),
            .lcout(chary_if_generate_plus_mult1_un68_sum_0_0_0_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2TEJF4_0_4_LC_5_4_2.C_ON=1'b0;
    defparam beamY_RNI2TEJF4_0_4_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2TEJF4_0_4_LC_5_4_2.LUT_INIT=16'b0101010101100110;
    LogicCell40 beamY_RNI2TEJF4_0_4_LC_5_4_2 (
            .in0(N__10046),
            .in1(N__9846),
            .in2(_gnd_net_),
            .in3(N__9256),
            .lcout(chary_if_generate_plus_mult1_un61_sum_0_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_0_3_LC_5_4_3.C_ON=1'b0;
    defparam beamY_RNIHUG2_0_3_LC_5_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_0_3_LC_5_4_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNIHUG2_0_3_LC_5_4_3 (
            .in0(_gnd_net_),
            .in1(N__10662),
            .in2(_gnd_net_),
            .in3(N__12247),
            .lcout(un5_visibley_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ53PA3_4_LC_5_4_4.C_ON=1'b0;
    defparam beamY_RNIQ53PA3_4_LC_5_4_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ53PA3_4_LC_5_4_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 beamY_RNIQ53PA3_4_LC_5_4_4 (
            .in0(_gnd_net_),
            .in1(N__9845),
            .in2(_gnd_net_),
            .in3(N__9255),
            .lcout(chary_if_generate_plus_mult1_un61_sum_c5),
            .ltout(chary_if_generate_plus_mult1_un61_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIUAPPF4_3_LC_5_4_5.C_ON=1'b0;
    defparam beamY_RNIUAPPF4_3_LC_5_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIUAPPF4_3_LC_5_4_5.LUT_INIT=16'b0010101110110010;
    LogicCell40 beamY_RNIUAPPF4_3_LC_5_4_5 (
            .in0(N__8443),
            .in1(N__9770),
            .in2(N__8437),
            .in3(N__10047),
            .lcout(chary_if_generate_plus_mult1_un68_sum_c4_0),
            .ltout(chary_if_generate_plus_mult1_un68_sum_c4_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKP1Q9A_5_LC_5_4_6.C_ON=1'b0;
    defparam beamY_RNIKP1Q9A_5_LC_5_4_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIKP1Q9A_5_LC_5_4_6.LUT_INIT=16'b1011001001110001;
    LogicCell40 beamY_RNIKP1Q9A_5_LC_5_4_6 (
            .in0(N__8401),
            .in1(N__8433),
            .in2(N__8425),
            .in3(N__9923),
            .lcout(),
            .ltout(g1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBLQCVR_2_LC_5_4_7.C_ON=1'b0;
    defparam beamY_RNIBLQCVR_2_LC_5_4_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIBLQCVR_2_LC_5_4_7.LUT_INIT=16'b0000000001101001;
    LogicCell40 beamY_RNIBLQCVR_2_LC_5_4_7 (
            .in0(N__8422),
            .in1(N__9322),
            .in2(N__8416),
            .in3(N__12248),
            .lcout(g2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIV142B4_3_LC_5_5_0.C_ON=1'b0;
    defparam beamY_RNIV142B4_3_LC_5_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIV142B4_3_LC_5_5_0.LUT_INIT=16'b1111111101101001;
    LogicCell40 beamY_RNIV142B4_3_LC_5_5_0 (
            .in0(N__9910),
            .in1(N__9348),
            .in2(N__9297),
            .in3(N__10642),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un75_sum_c5_N_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICECPQ8_4_LC_5_5_1.C_ON=1'b0;
    defparam beamY_RNICECPQ8_4_LC_5_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNICECPQ8_4_LC_5_5_1.LUT_INIT=16'b1011100011100010;
    LogicCell40 beamY_RNICECPQ8_4_LC_5_5_1 (
            .in0(N__8413),
            .in1(N__9190),
            .in2(N__8404),
            .in3(N__8647),
            .lcout(chary_if_generate_plus_mult1_un75_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFJKLC_0_5_LC_5_5_2.C_ON=1'b0;
    defparam beamY_RNIFJKLC_0_5_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIFJKLC_0_5_LC_5_5_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIFJKLC_0_5_LC_5_5_2 (
            .in0(N__9720),
            .in1(N__10085),
            .in2(N__9638),
            .in3(N__9545),
            .lcout(g0_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKHPCA1_5_LC_5_5_3.C_ON=1'b0;
    defparam beamY_RNIKHPCA1_5_LC_5_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIKHPCA1_5_LC_5_5_3.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIKHPCA1_5_LC_5_5_3 (
            .in0(N__10086),
            .in1(N__9630),
            .in2(N__8395),
            .in3(N__9911),
            .lcout(chary_if_generate_plus_mult1_un61_sum_1_0_1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI44RHC_5_LC_5_5_4.C_ON=1'b0;
    defparam beamY_RNI44RHC_5_LC_5_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI44RHC_5_LC_5_5_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNI44RHC_5_LC_5_5_4 (
            .in0(N__9626),
            .in1(N__10084),
            .in2(_gnd_net_),
            .in3(N__9542),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNINITP61_5_LC_5_5_5.C_ON=1'b0;
    defparam beamY_RNINITP61_5_LC_5_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNINITP61_5_LC_5_5_5.LUT_INIT=16'b1000111011010100;
    LogicCell40 beamY_RNINITP61_5_LC_5_5_5 (
            .in0(N__9544),
            .in1(N__10135),
            .in2(N__9739),
            .in3(N__9909),
            .lcout(),
            .ltout(beamY_RNINITP61Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITFRN03_5_LC_5_5_6.C_ON=1'b0;
    defparam beamY_RNITFRN03_5_LC_5_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNITFRN03_5_LC_5_5_6.LUT_INIT=16'b1111001111000000;
    LogicCell40 beamY_RNITFRN03_5_LC_5_5_6 (
            .in0(_gnd_net_),
            .in1(N__9137),
            .in2(N__8488),
            .in3(N__8485),
            .lcout(beamY_RNITFRN03Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNINITP61_1_5_LC_5_5_7.C_ON=1'b0;
    defparam beamY_RNINITP61_1_5_LC_5_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNINITP61_1_5_LC_5_5_7.LUT_INIT=16'b0111000100101011;
    LogicCell40 beamY_RNINITP61_1_5_LC_5_5_7 (
            .in0(N__9543),
            .in1(N__10134),
            .in2(N__9738),
            .in3(N__9908),
            .lcout(beamY_RNINITP61_1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIIIGJ2_0_9_LC_5_6_0.C_ON=1'b0;
    defparam beamY_RNIIIGJ2_0_9_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIIIGJ2_0_9_LC_5_6_0.LUT_INIT=16'b0100101001011110;
    LogicCell40 beamY_RNIIIGJ2_0_9_LC_5_6_0 (
            .in0(N__8478),
            .in1(N__9403),
            .in2(N__12809),
            .in3(N__9803),
            .lcout(chary_if_generate_plus_mult1_un47_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIIIGJ2_9_LC_5_6_1.C_ON=1'b0;
    defparam beamY_RNIIIGJ2_9_LC_5_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIIIGJ2_9_LC_5_6_1.LUT_INIT=16'b1001110000111001;
    LogicCell40 beamY_RNIIIGJ2_9_LC_5_6_1 (
            .in0(N__12792),
            .in1(N__8479),
            .in2(N__9816),
            .in3(N__9427),
            .lcout(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0),
            .ltout(chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI14TP8_7_LC_5_6_2.C_ON=1'b0;
    defparam beamY_RNI14TP8_7_LC_5_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI14TP8_7_LC_5_6_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNI14TP8_7_LC_5_6_2 (
            .in0(N__8701),
            .in1(N__8467),
            .in2(N__8470),
            .in3(N__8458),
            .lcout(chary_if_generate_plus_mult1_un54_sum_axbxc5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITKMQ1_9_LC_5_6_3.C_ON=1'b0;
    defparam beamY_RNITKMQ1_9_LC_5_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNITKMQ1_9_LC_5_6_3.LUT_INIT=16'b1010101010011001;
    LogicCell40 beamY_RNITKMQ1_9_LC_5_6_3 (
            .in0(N__9808),
            .in1(N__12670),
            .in2(_gnd_net_),
            .in3(N__12584),
            .lcout(chary_if_generate_plus_mult1_un47_sum_axbxc5_2),
            .ltout(chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIB65I6_7_LC_5_6_4.C_ON=1'b0;
    defparam beamY_RNIB65I6_7_LC_5_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIB65I6_7_LC_5_6_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIB65I6_7_LC_5_6_4 (
            .in0(N__8700),
            .in1(N__8457),
            .in2(N__8461),
            .in3(N__9404),
            .lcout(chary_if_generate_plus_mult1_un54_sum_axb3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITURI3_7_LC_5_6_5.C_ON=1'b0;
    defparam beamY_RNITURI3_7_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNITURI3_7_LC_5_6_5.LUT_INIT=16'b1010010110010110;
    LogicCell40 beamY_RNITURI3_7_LC_5_6_5 (
            .in0(N__8455),
            .in1(N__12666),
            .in2(N__9815),
            .in3(N__12582),
            .lcout(beamY_RNITURI3Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITURI3_0_7_LC_5_6_6.C_ON=1'b0;
    defparam beamY_RNITURI3_0_7_LC_5_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNITURI3_0_7_LC_5_6_6.LUT_INIT=16'b0011011011001001;
    LogicCell40 beamY_RNITURI3_0_7_LC_5_6_6 (
            .in0(N__12583),
            .in1(N__8456),
            .in2(N__12686),
            .in3(N__9804),
            .lcout(),
            .ltout(beamY_RNITURI3_0Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNICG8P9_7_LC_5_6_7.C_ON=1'b0;
    defparam beamY_RNICG8P9_7_LC_5_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNICG8P9_7_LC_5_6_7.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNICG8P9_7_LC_5_6_7 (
            .in0(_gnd_net_),
            .in1(N__8699),
            .in2(N__8689),
            .in3(N__8686),
            .lcout(beamY_RNICG8P9Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un15_beamy_2_LC_5_7_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un15_beamy_2_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un15_beamy_2_LC_5_7_0.LUT_INIT=16'b0000000000000001;
    LogicCell40 un114_pixel_1_0_3__un15_beamy_2_LC_5_7_0 (
            .in0(N__8554),
            .in1(N__8680),
            .in2(N__10237),
            .in3(N__8674),
            .lcout(un114_pixel_1_0_3__un15_beamyZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un3_beamx_2_LC_5_7_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un3_beamx_2_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un3_beamx_2_LC_5_7_1.LUT_INIT=16'b0000000000110011;
    LogicCell40 un114_pixel_1_0_3__un3_beamx_2_LC_5_7_1 (
            .in0(_gnd_net_),
            .in1(N__10746),
            .in2(_gnd_net_),
            .in3(N__10281),
            .lcout(un1_beamx_2),
            .ltout(un1_beamx_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un15_beamy_LC_5_7_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un15_beamy_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un15_beamy_LC_5_7_2.LUT_INIT=16'b0100110000001100;
    LogicCell40 un114_pixel_1_0_3__un15_beamy_LC_5_7_2 (
            .in0(N__8755),
            .in1(N__8668),
            .in2(N__8662),
            .in3(N__10322),
            .lcout(un15_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un5_beamx_3_LC_5_7_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un5_beamx_3_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un5_beamx_3_LC_5_7_5.LUT_INIT=16'b0000000001000100;
    LogicCell40 un114_pixel_1_0_3__un5_beamx_3_LC_5_7_5 (
            .in0(N__14634),
            .in1(N__10667),
            .in2(_gnd_net_),
            .in3(N__12253),
            .lcout(un114_pixel_1_0_3__un5_beamxZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_1_3_LC_5_7_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_1_3_LC_5_7_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_1_3_LC_5_7_6.LUT_INIT=16'b0000000000010011;
    LogicCell40 un114_pixel_1_0_3__g0_1_3_LC_5_7_6 (
            .in0(N__12254),
            .in1(N__10668),
            .in2(N__15016),
            .in3(N__8646),
            .lcout(un114_pixel_1_0_3__g0_1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un18_beamylto9_2_LC_5_8_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un18_beamylto9_2_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un18_beamylto9_2_LC_5_8_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_1_0_3__un18_beamylto9_2_LC_5_8_0 (
            .in0(N__10273),
            .in1(N__10312),
            .in2(N__10747),
            .in3(N__10364),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un18_beamylto9Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un18_beamylto9_LC_5_8_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un18_beamylto9_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un18_beamylto9_LC_5_8_1.LUT_INIT=16'b1101000011000000;
    LogicCell40 un114_pixel_1_0_3__un18_beamylto9_LC_5_8_1 (
            .in0(N__10188),
            .in1(N__10397),
            .in2(N__8557),
            .in3(N__10448),
            .lcout(un18_beamylt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_1_LC_5_8_3.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_1_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_1_LC_5_8_3.LUT_INIT=16'b0111000000110101;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_1_LC_5_8_3 (
            .in0(N__12251),
            .in1(N__8545),
            .in2(N__8749),
            .in3(N__10663),
            .lcout(row_1_if_generate_plus_mult1_un82_sum_ac0_7_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un13_beamylto6_LC_5_8_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un13_beamylto6_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un13_beamylto6_LC_5_8_4.LUT_INIT=16'b0011001100010011;
    LogicCell40 un114_pixel_1_0_3__un13_beamylto6_LC_5_8_4 (
            .in0(N__10449),
            .in1(N__10365),
            .in2(N__10411),
            .in3(N__10189),
            .lcout(un13_beamylt7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_LC_5_8_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_LC_5_8_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_axb4_LC_5_8_6.LUT_INIT=16'b1001011001101001;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_axb4_LC_5_8_6 (
            .in0(N__12438),
            .in1(N__8736),
            .in2(N__12465),
            .in3(N__12406),
            .lcout(),
            .ltout(row_1_if_generate_plus_mult1_un82_sum_axb4_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_5_8_7.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_5_8_7.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_5_8_7.LUT_INIT=16'b0100111101000100;
    LogicCell40 row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_5_8_7 (
            .in0(N__8748),
            .in1(N__8737),
            .in2(N__8725),
            .in3(N__8722),
            .lcout(row_1_if_generate_plus_mult1_un82_sum_c5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_5_9_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_5_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_5_9_0 (
            .in0(_gnd_net_),
            .in1(N__10550),
            .in2(N__12024),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_5_9_1.C_ON=1'b1;
    defparam beamX_2_LC_5_9_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_5_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(N__10518),
            .in2(_gnd_net_),
            .in3(N__8716),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__11874),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_5_9_2.C_ON=1'b1;
    defparam beamX_3_LC_5_9_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_5_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_5_9_2 (
            .in0(_gnd_net_),
            .in1(N__10486),
            .in2(_gnd_net_),
            .in3(N__8713),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__11874),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_5_9_3.C_ON=1'b1;
    defparam beamX_4_LC_5_9_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_5_9_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_5_9_3 (
            .in0(N__11040),
            .in1(N__10451),
            .in2(_gnd_net_),
            .in3(N__8710),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__11874),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_5_9_4.C_ON=1'b1;
    defparam beamX_5_LC_5_9_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_5_9_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_5_9_4 (
            .in0(_gnd_net_),
            .in1(N__10414),
            .in2(_gnd_net_),
            .in3(N__8707),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__11874),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_5_9_5.C_ON=1'b1;
    defparam beamX_6_LC_5_9_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_5_9_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_5_9_5 (
            .in0(_gnd_net_),
            .in1(N__10367),
            .in2(_gnd_net_),
            .in3(N__8704),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__11874),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_5_9_6.C_ON=1'b1;
    defparam beamX_7_LC_5_9_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_5_9_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_5_9_6 (
            .in0(_gnd_net_),
            .in1(N__10321),
            .in2(_gnd_net_),
            .in3(N__8779),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__11874),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_5_9_7.C_ON=1'b1;
    defparam beamX_8_LC_5_9_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_5_9_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_5_9_7 (
            .in0(_gnd_net_),
            .in1(N__10277),
            .in2(_gnd_net_),
            .in3(N__8776),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__11874),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_5_10_0.C_ON=1'b1;
    defparam beamX_9_LC_5_10_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_5_10_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_5_10_0 (
            .in0(_gnd_net_),
            .in1(N__10742),
            .in2(_gnd_net_),
            .in3(N__8773),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__11879),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_5_10_1.C_ON=1'b0;
    defparam beamX_10_LC_5_10_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_5_10_1.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamX_10_LC_5_10_1 (
            .in0(N__10231),
            .in1(N__11042),
            .in2(_gnd_net_),
            .in3(N__8770),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11879),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8V_LC_5_10_3.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8V_LC_5_10_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8V_LC_5_10_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8V_LC_5_10_3 (
            .in0(_gnd_net_),
            .in1(N__10174),
            .in2(_gnd_net_),
            .in3(N__10175),
            .lcout(charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8VZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_5_10_4.C_ON=1'b0;
    defparam beamX_1_LC_5_10_4.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_5_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamX_1_LC_5_10_4 (
            .in0(_gnd_net_),
            .in1(N__10551),
            .in2(_gnd_net_),
            .in3(N__12002),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11879),
            .ce(),
            .sr(_gnd_net_));
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_2_LC_5_10_6.C_ON=1'b0;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_2_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_2_LC_5_10_6.LUT_INIT=16'b0010110101001011;
    LogicCell40 row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_2_LC_5_10_6 (
            .in0(N__12723),
            .in1(N__9784),
            .in2(N__8767),
            .in3(N__9592),
            .lcout(row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__N_204_0_i_LC_5_11_0.C_ON=1'b1;
    defparam un114_pixel_1_0_3__N_204_0_i_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__N_204_0_i_LC_5_11_0.LUT_INIT=16'b0000111111111111;
    LogicCell40 un114_pixel_1_0_3__N_204_0_i_LC_5_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16155),
            .in3(N__12937),
            .lcout(N_204_0_i),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(charx_if_generate_plus_mult1_un19_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_LUT4_0_LC_5_11_1.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_LUT4_0_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_LUT4_0_LC_5_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_LUT4_0_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8758),
            .lcout(charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_5_11_4.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_0_LC_5_11_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_0_LC_5_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13872),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_5_11_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_5_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_0_LC_5_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_0_LC_5_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11649),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam nCS1_1_RNO_0_LC_5_13_2.C_ON=1'b0;
    defparam nCS1_1_RNO_0_LC_5_13_2.SEQ_MODE=4'b0000;
    defparam nCS1_1_RNO_0_LC_5_13_2.LUT_INIT=16'b1000100011001000;
    LogicCell40 nCS1_1_RNO_0_LC_5_13_2 (
            .in0(N__9024),
            .in1(N__8893),
            .in2(N__8940),
            .in3(N__9000),
            .lcout(nCS1_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_5_LC_5_13_4.C_ON=1'b0;
    defparam counter_5_LC_5_13_4.SEQ_MODE=4'b1000;
    defparam counter_5_LC_5_13_4.LUT_INIT=16'b1000100000001100;
    LogicCell40 counter_5_LC_5_13_4 (
            .in0(N__8968),
            .in1(N__9031),
            .in2(N__8860),
            .in3(N__8898),
            .lcout(counterZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14327),
            .ce(),
            .sr(_gnd_net_));
    defparam slaveselect_LC_5_13_5.C_ON=1'b0;
    defparam slaveselect_LC_5_13_5.SEQ_MODE=4'b1000;
    defparam slaveselect_LC_5_13_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 slaveselect_LC_5_13_5 (
            .in0(N__8894),
            .in1(N__8854),
            .in2(_gnd_net_),
            .in3(N__8966),
            .lcout(slaveselectZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14327),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_RNIQHKU_5_LC_5_13_6.C_ON=1'b0;
    defparam counter_RNIQHKU_5_LC_5_13_6.SEQ_MODE=4'b0000;
    defparam counter_RNIQHKU_5_LC_5_13_6.LUT_INIT=16'b1100100011001100;
    LogicCell40 counter_RNIQHKU_5_LC_5_13_6 (
            .in0(N__9025),
            .in1(N__8899),
            .in2(N__8941),
            .in3(N__9001),
            .lcout(un1_slaveselect_1_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam counter_4_LC_5_13_7.C_ON=1'b0;
    defparam counter_4_LC_5_13_7.SEQ_MODE=4'b1000;
    defparam counter_4_LC_5_13_7.LUT_INIT=16'b1100010100000000;
    LogicCell40 counter_4_LC_5_13_7 (
            .in0(N__8853),
            .in1(N__8967),
            .in2(N__8909),
            .in3(N__8947),
            .lcout(counterZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14327),
            .ce(),
            .sr(_gnd_net_));
    defparam nCS1_1_LC_5_14_5.C_ON=1'b0;
    defparam nCS1_1_LC_5_14_5.SEQ_MODE=4'b1001;
    defparam nCS1_1_LC_5_14_5.LUT_INIT=16'b1000100010111011;
    LogicCell40 nCS1_1_LC_5_14_5 (
            .in0(N__8802),
            .in1(N__8908),
            .in2(_gnd_net_),
            .in3(N__8859),
            .lcout(nCS1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14328),
            .ce(),
            .sr(N__8791));
    defparam un114_pixel_1_0_3__g0_8_LC_6_3_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_8_LC_6_3_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_8_LC_6_3_0.LUT_INIT=16'b1000010000010010;
    LogicCell40 un114_pixel_1_0_3__g0_8_LC_6_3_0 (
            .in0(N__9360),
            .in1(N__9088),
            .in2(N__9112),
            .in3(N__12250),
            .lcout(font_un28_pixel_0_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2TEJF4_4_LC_6_3_2.C_ON=1'b0;
    defparam beamY_RNI2TEJF4_4_LC_6_3_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2TEJF4_4_LC_6_3_2.LUT_INIT=16'b0101010101100110;
    LogicCell40 beamY_RNI2TEJF4_4_LC_6_3_2 (
            .in0(N__10043),
            .in1(N__9857),
            .in2(_gnd_net_),
            .in3(N__9254),
            .lcout(beamY_RNI2TEJF4Z0Z_4),
            .ltout(beamY_RNI2TEJF4Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_8_1_LC_6_3_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_8_1_LC_6_3_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_8_1_LC_6_3_3.LUT_INIT=16'b0111111010000001;
    LogicCell40 un114_pixel_1_0_3__g0_8_1_LC_6_3_3 (
            .in0(N__9221),
            .in1(N__9163),
            .in2(N__9115),
            .in3(N__10664),
            .lcout(un114_pixel_1_0_3__g0_8Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKHPCA1_0_4_LC_6_3_4.C_ON=1'b0;
    defparam beamY_RNIKHPCA1_0_4_LC_6_3_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIKHPCA1_0_4_LC_6_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNIKHPCA1_0_4_LC_6_3_4 (
            .in0(N__9769),
            .in1(N__9295),
            .in2(_gnd_net_),
            .in3(N__9932),
            .lcout(chary_if_generate_plus_mult1_un61_sum_0_3),
            .ltout(chary_if_generate_plus_mult1_un61_sum_0_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_10_LC_6_3_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_10_LC_6_3_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_10_LC_6_3_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un114_pixel_1_0_3__g0_10_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(N__10044),
            .in2(N__9103),
            .in3(N__9359),
            .lcout(),
            .ltout(un114_pixel_1_0_3__g0_1Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_3_0_LC_6_3_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_3_0_LC_6_3_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_3_0_LC_6_3_6.LUT_INIT=16'b0001111011100001;
    LogicCell40 un114_pixel_1_0_3__g0_3_0_LC_6_3_6 (
            .in0(N__9259),
            .in1(N__9858),
            .in2(N__9100),
            .in3(N__9325),
            .lcout(),
            .ltout(un114_pixel_1_0_3__g0_3Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_9_LC_6_3_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_9_LC_6_3_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_9_LC_6_3_7.LUT_INIT=16'b1000011111100001;
    LogicCell40 un114_pixel_1_0_3__g0_9_LC_6_3_7 (
            .in0(N__9097),
            .in1(N__9186),
            .in2(N__9091),
            .in3(N__9162),
            .lcout(chary_if_generate_plus_mult1_un75_sum_i_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_6_LC_6_4_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_6_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_6_LC_6_4_0.LUT_INIT=16'b0011110001101001;
    LogicCell40 un114_pixel_1_0_3__g0_6_LC_6_4_0 (
            .in0(N__9855),
            .in1(N__10035),
            .in2(N__9952),
            .in3(N__9258),
            .lcout(),
            .ltout(un114_pixel_1_0_3__g0Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_5_LC_6_4_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_5_LC_6_4_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_5_LC_6_4_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un114_pixel_1_0_3__g0_5_LC_6_4_1 (
            .in0(_gnd_net_),
            .in1(N__9082),
            .in2(N__9070),
            .in3(N__9323),
            .lcout(),
            .ltout(un114_pixel_1_0_3__g0Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_0_1_LC_6_4_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_0_1_LC_6_4_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_0_1_LC_6_4_2.LUT_INIT=16'b1101101101111110;
    LogicCell40 un114_pixel_1_0_3__g0_0_1_LC_6_4_2 (
            .in0(N__9067),
            .in1(N__9061),
            .in2(N__9055),
            .in3(N__10665),
            .lcout(un114_pixel_1_0_3__N_5_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIH9THAD_4_LC_6_4_3.C_ON=1'b0;
    defparam beamY_RNIH9THAD_4_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIH9THAD_4_LC_6_4_3.LUT_INIT=16'b0111111010000001;
    LogicCell40 beamY_RNIH9THAD_4_LC_6_4_3 (
            .in0(N__9184),
            .in1(N__9159),
            .in2(N__9226),
            .in3(N__9357),
            .lcout(beamY_RNIH9THADZ0Z_4),
            .ltout(beamY_RNIH9THADZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHHB5F01_4_LC_6_4_4.C_ON=1'b0;
    defparam beamY_RNIHHB5F01_4_LC_6_4_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIHHB5F01_4_LC_6_4_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIHHB5F01_4_LC_6_4_4 (
            .in0(N__9324),
            .in1(N__9196),
            .in2(N__9301),
            .in3(N__9161),
            .lcout(beamY_RNIHHB5F01Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI3SPGT1_4_LC_6_4_5.C_ON=1'b0;
    defparam beamY_RNI3SPGT1_4_LC_6_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI3SPGT1_4_LC_6_4_5.LUT_INIT=16'b0010000001000000;
    LogicCell40 beamY_RNI3SPGT1_4_LC_6_4_5 (
            .in0(N__9139),
            .in1(N__9282),
            .in2(N__9781),
            .in3(N__9906),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_7_d),
            .ltout(chary_if_generate_plus_mult1_un61_sum_ac0_7_d_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIME80Q5_4_LC_6_4_6.C_ON=1'b0;
    defparam beamY_RNIME80Q5_4_LC_6_4_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIME80Q5_4_LC_6_4_6.LUT_INIT=16'b0011011011001001;
    LogicCell40 beamY_RNIME80Q5_4_LC_6_4_6 (
            .in0(N__9856),
            .in1(N__9222),
            .in2(N__9199),
            .in3(N__10034),
            .lcout(chary_if_generate_plus_mult1_un68_sum_axb4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKP1Q9A_0_5_LC_6_4_7.C_ON=1'b0;
    defparam beamY_RNIKP1Q9A_0_5_LC_6_4_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIKP1Q9A_0_5_LC_6_4_7.LUT_INIT=16'b0001100010000001;
    LogicCell40 beamY_RNIKP1Q9A_0_5_LC_6_4_7 (
            .in0(N__9185),
            .in1(N__9160),
            .in2(N__9604),
            .in3(N__9907),
            .lcout(g1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFA04J_5_LC_6_5_0.C_ON=1'b0;
    defparam beamY_RNIFA04J_5_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIFA04J_5_LC_6_5_0.LUT_INIT=16'b1001011001101001;
    LogicCell40 beamY_RNIFA04J_5_LC_6_5_0 (
            .in0(N__9539),
            .in1(N__9479),
            .in2(N__9639),
            .in3(N__10083),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGS0LB_5_LC_6_5_1.C_ON=1'b0;
    defparam beamY_RNIGS0LB_5_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIGS0LB_5_LC_6_5_1.LUT_INIT=16'b1101010011110100;
    LogicCell40 beamY_RNIGS0LB_5_LC_6_5_1 (
            .in0(N__10082),
            .in1(N__9538),
            .in2(N__10111),
            .in3(N__9450),
            .lcout(beamY_RNIGS0LBZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNINITP61_0_5_LC_6_5_2.C_ON=1'b0;
    defparam beamY_RNINITP61_0_5_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNINITP61_0_5_LC_6_5_2.LUT_INIT=16'b0111000100101011;
    LogicCell40 beamY_RNINITP61_0_5_LC_6_5_2 (
            .in0(N__9541),
            .in1(N__10138),
            .in2(N__9760),
            .in3(N__9924),
            .lcout(),
            .ltout(g0_0_x2_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVC6VP1_3_LC_6_5_3.C_ON=1'b0;
    defparam beamY_RNIVC6VP1_3_LC_6_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIVC6VP1_3_LC_6_5_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamY_RNIVC6VP1_3_LC_6_5_3 (
            .in0(_gnd_net_),
            .in1(N__9138),
            .in2(N__9118),
            .in3(N__10658),
            .lcout(g0_0_x2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIC02EA1_2_LC_6_5_4.C_ON=1'b0;
    defparam beamY_RNIC02EA1_2_LC_6_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIC02EA1_2_LC_6_5_4.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIC02EA1_2_LC_6_5_4 (
            .in0(N__9721),
            .in1(N__9823),
            .in2(N__9931),
            .in3(N__12249),
            .lcout(g0_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIARUFB_5_LC_6_5_5.C_ON=1'b0;
    defparam beamY_RNIARUFB_5_LC_6_5_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIARUFB_5_LC_6_5_5.LUT_INIT=16'b0010001010101010;
    LogicCell40 beamY_RNIARUFB_5_LC_6_5_5 (
            .in0(N__10109),
            .in1(N__10081),
            .in2(_gnd_net_),
            .in3(N__9451),
            .lcout(),
            .ltout(beamY_RNIARUFBZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5U4NT_5_LC_6_5_6.C_ON=1'b0;
    defparam beamY_RNI5U4NT_5_LC_6_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI5U4NT_5_LC_6_5_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNI5U4NT_5_LC_6_5_6 (
            .in0(_gnd_net_),
            .in1(N__9478),
            .in2(N__9943),
            .in3(N__9940),
            .lcout(chary_if_generate_plus_mult1_un54_sum_c5),
            .ltout(chary_if_generate_plus_mult1_un54_sum_c5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN998D1_5_LC_6_5_7.C_ON=1'b0;
    defparam beamY_RNIN998D1_5_LC_6_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIN998D1_5_LC_6_5_7.LUT_INIT=16'b0100000110101010;
    LogicCell40 beamY_RNIN998D1_5_LC_6_5_7 (
            .in0(N__9480),
            .in1(N__10136),
            .in2(N__9862),
            .in3(N__9540),
            .lcout(chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI44RHC_0_5_LC_6_6_1.C_ON=1'b0;
    defparam beamY_RNI44RHC_0_5_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI44RHC_0_5_LC_6_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_RNI44RHC_0_5_LC_6_6_1 (
            .in0(N__9588),
            .in1(N__9634),
            .in2(_gnd_net_),
            .in3(N__10089),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axb3_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2MTA1_9_LC_6_6_2.C_ON=1'b0;
    defparam beamY_RNI2MTA1_9_LC_6_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2MTA1_9_LC_6_6_2.LUT_INIT=16'b0110011010011001;
    LogicCell40 beamY_RNI2MTA1_9_LC_6_6_2 (
            .in0(N__9817),
            .in1(N__9458),
            .in2(_gnd_net_),
            .in3(N__12791),
            .lcout(beamY_RNI2MTA1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIFJKLC_5_LC_6_6_4.C_ON=1'b0;
    defparam beamY_RNIFJKLC_5_LC_6_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIFJKLC_5_LC_6_6_4.LUT_INIT=16'b0110100110010110;
    LogicCell40 beamY_RNIFJKLC_5_LC_6_6_4 (
            .in0(N__10090),
            .in1(N__9780),
            .in2(N__9640),
            .in3(N__9589),
            .lcout(g0_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPC8SG_5_LC_6_6_6.C_ON=1'b0;
    defparam beamY_RNIPC8SG_5_LC_6_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIPC8SG_5_LC_6_6_6.LUT_INIT=16'b1100000011101010;
    LogicCell40 beamY_RNIPC8SG_5_LC_6_6_6 (
            .in0(N__10087),
            .in1(N__9587),
            .in2(N__9484),
            .in3(N__9459),
            .lcout(),
            .ltout(chary_if_generate_plus_mult1_un54_sum_c4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI8NBQ41_5_LC_6_6_7.C_ON=1'b0;
    defparam beamY_RNI8NBQ41_5_LC_6_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNI8NBQ41_5_LC_6_6_7.LUT_INIT=16'b1010100101101010;
    LogicCell40 beamY_RNI8NBQ41_5_LC_6_6_7 (
            .in0(N__10137),
            .in1(N__10110),
            .in2(N__10093),
            .in3(N__10088),
            .lcout(chary_if_generate_plus_mult1_un61_sum_axbxc5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un3_beamx_LC_6_7_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un3_beamx_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un3_beamx_LC_6_7_2.LUT_INIT=16'b0000000000001000;
    LogicCell40 un114_pixel_1_0_3__un3_beamx_LC_6_7_2 (
            .in0(N__10198),
            .in1(N__9996),
            .in2(N__10329),
            .in3(N__10412),
            .lcout(un3_beamx_0),
            .ltout(un3_beamx_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_6_7_3.C_ON=1'b0;
    defparam beamY_0_LC_6_7_3.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_6_7_3.LUT_INIT=16'b0000111100110000;
    LogicCell40 beamY_0_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(N__10970),
            .in2(N__10000),
            .in3(N__14641),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11881),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJPPPPD1_3_LC_6_7_4.C_ON=1'b0;
    defparam beamY_RNIJPPPPD1_3_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIJPPPPD1_3_LC_6_7_4.LUT_INIT=16'b0011110010010110;
    LogicCell40 beamY_RNIJPPPPD1_3_LC_6_7_4 (
            .in0(N__12291),
            .in1(N__10666),
            .in2(N__10690),
            .in3(N__12252),
            .lcout(chary_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSyncZ0_LC_6_7_6.C_ON=1'b0;
    defparam HSyncZ0_LC_6_7_6.SEQ_MODE=4'b1000;
    defparam HSyncZ0_LC_6_7_6.LUT_INIT=16'b1111111111111011;
    LogicCell40 HSyncZ0_LC_6_7_6 (
            .in0(N__10236),
            .in1(N__9997),
            .in2(N__10330),
            .in3(N__10243),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11881),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_6_8_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_6_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_6_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15093),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_6_8_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_6_8_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_6_8_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_6_8_1 (
            .in0(_gnd_net_),
            .in1(N__10144),
            .in2(_gnd_net_),
            .in3(N__9973),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HL_LC_6_8_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HL_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HL_LC_6_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HL_LC_6_8_2 (
            .in0(_gnd_net_),
            .in1(N__16364),
            .in2(N__10153),
            .in3(N__9970),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HLZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_c_RNIMVPQ1_LC_6_8_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_c_RNIMVPQ1_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_3_c_RNIMVPQ1_LC_6_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_3_c_RNIMVPQ1_LC_6_8_3 (
            .in0(N__11229),
            .in1(N__10180),
            .in2(N__9967),
            .in3(N__9955),
            .lcout(charx_if_generate_plus_mult1_un33_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un26_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un26_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_6_8_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_6_8_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_6_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10246),
            .lcout(charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un1_beamxlto6_LC_6_8_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un1_beamxlto6_LC_6_8_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un1_beamxlto6_LC_6_8_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_1_0_3__un1_beamxlto6_LC_6_8_6 (
            .in0(N__10413),
            .in1(N__10452),
            .in2(N__10492),
            .in3(N__10368),
            .lcout(un1_beamxlt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un3_beamx_5_LC_6_9_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un3_beamx_5_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un3_beamx_5_LC_6_9_0.LUT_INIT=16'b0001000000000000;
    LogicCell40 un114_pixel_1_0_3__un3_beamx_5_LC_6_9_0 (
            .in0(N__10549),
            .in1(N__10517),
            .in2(N__10235),
            .in3(N__10450),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un3_beamxZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un3_beamx_7_LC_6_9_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un3_beamx_7_LC_6_9_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un3_beamx_7_LC_6_9_1.LUT_INIT=16'b0000000000010000;
    LogicCell40 un114_pixel_1_0_3__un3_beamx_7_LC_6_9_1 (
            .in0(N__10485),
            .in1(N__10366),
            .in2(N__10201),
            .in3(N__11989),
            .lcout(un114_pixel_1_0_3__un3_beamxZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_4_0_15__un13_beamylto3_LC_6_9_3.C_ON=1'b0;
    defparam un114_pixel_4_0_15__un13_beamylto3_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_4_0_15__un13_beamylto3_LC_6_9_3.LUT_INIT=16'b0000011100001111;
    LogicCell40 un114_pixel_4_0_15__un13_beamylto3_LC_6_9_3 (
            .in0(N__10516),
            .in1(N__10548),
            .in2(N__10491),
            .in3(N__11988),
            .lcout(un18_beamylt4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_6_9_4.C_ON=1'b0;
    defparam beamX_0_LC_6_9_4.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_6_9_4.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamX_0_LC_6_9_4 (
            .in0(N__11990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11041),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11876),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKF_LC_6_9_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKF_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKF_LC_6_9_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKF_LC_6_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10179),
            .lcout(charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKFZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_N_575_i_LC_6_9_6.C_ON=1'b0;
    defparam column_1_N_575_i_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam column_1_N_575_i_LC_6_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_N_575_i_LC_6_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11645),
            .lcout(N_575_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_6_9_7.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_6_9_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_1_LC_6_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_1_LC_6_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16156),
            .lcout(charx_if_generate_plus_mult1_un19_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_LC_6_10_0.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_LC_6_10_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_LC_6_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_cry_0_c_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12003),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(un5_visiblex_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_6_10_1.C_ON=1'b1;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_6_10_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_0_c_RNIHKT1_LC_6_10_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_0_c_RNIHKT1_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10552),
            .in3(N__10522),
            .lcout(charx_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_0),
            .carryout(un5_visiblex_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_6_10_2.C_ON=1'b1;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_6_10_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_LC_6_10_2.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_LC_6_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10519),
            .in3(N__10495),
            .lcout(charx_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_1),
            .carryout(un5_visiblex_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_6_10_3.C_ON=1'b1;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_6_10_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_LC_6_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_LC_6_10_3 (
            .in0(_gnd_net_),
            .in1(N__16394),
            .in2(N__10490),
            .in3(N__10456),
            .lcout(chessboardpixel_un152_pixel_24),
            .ltout(),
            .carryin(un5_visiblex_cry_2),
            .carryout(un5_visiblex_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_LC_6_10_4.C_ON=1'b1;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_LC_6_10_4.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_LC_6_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10453),
            .in3(N__10417),
            .lcout(charx_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_3),
            .carryout(un5_visiblex_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_LC_6_10_5.C_ON=1'b1;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_LC_6_10_5.LUT_INIT=16'b1010010101011010;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_LC_6_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10410),
            .in3(N__10372),
            .lcout(charx_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_4),
            .carryout(un5_visiblex_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_LC_6_10_6.C_ON=1'b1;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_6_10_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_LC_6_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_LC_6_10_6 (
            .in0(_gnd_net_),
            .in1(N__16395),
            .in2(N__10369),
            .in3(N__10333),
            .lcout(charx_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_5),
            .carryout(un5_visiblex_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_LC_6_10_7.C_ON=1'b1;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_6_10_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_LC_6_10_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_LC_6_10_7 (
            .in0(_gnd_net_),
            .in1(N__10311),
            .in2(_gnd_net_),
            .in3(N__10285),
            .lcout(charx_if_generate_plus_mult1_un33_sum),
            .ltout(),
            .carryin(un5_visiblex_cry_6),
            .carryout(un5_visiblex_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_LC_6_11_0.C_ON=1'b1;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_6_11_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_LC_6_11_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_LC_6_11_0 (
            .in0(_gnd_net_),
            .in1(N__16396),
            .in2(N__10282),
            .in3(N__10249),
            .lcout(charx_if_generate_plus_mult1_un26_sum),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(un5_visiblex_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_6_11_1.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_LC_6_11_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(N__10735),
            .in2(_gnd_net_),
            .in3(N__10714),
            .lcout(CO3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_4.C_ON=1'b0;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13876),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_3_bm_2_LC_7_3_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_3_bm_2_LC_7_3_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_3_bm_2_LC_7_3_0.LUT_INIT=16'b0000000011001111;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_3_bm_2_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__13417),
            .in2(N__16030),
            .in3(N__14750),
            .lcout(),
            .ltout(un116_pixel_3_bm_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_2_LC_7_3_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_2_LC_7_3_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_2_LC_7_3_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_3_ns_2_LC_7_3_1 (
            .in0(_gnd_net_),
            .in1(N__14949),
            .in2(N__10711),
            .in3(N__11662),
            .lcout(un116_pixel_3_ns_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_2_LC_7_3_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_2_LC_7_3_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_2_LC_7_3_2.LUT_INIT=16'b0000111001010000;
    LogicCell40 un114_pixel_1_0_3__g0_2_LC_7_3_2 (
            .in0(N__15814),
            .in1(N__10696),
            .in2(N__10708),
            .in3(N__15355),
            .lcout(N_345_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_16_LC_7_3_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_16_LC_7_3_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_16_LC_7_3_3.LUT_INIT=16'b0111001101010011;
    LogicCell40 un114_pixel_1_0_3__g0_16_LC_7_3_3 (
            .in0(N__15354),
            .in1(N__15813),
            .in2(N__14995),
            .in3(N__15585),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un116_pixel_4_ns_1_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_12_LC_7_3_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_12_LC_7_3_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_12_LC_7_3_4.LUT_INIT=16'b0100101010101110;
    LogicCell40 un114_pixel_1_0_3__g0_12_LC_7_3_4 (
            .in0(N__14950),
            .in1(N__14255),
            .in2(N__10699),
            .in3(N__16029),
            .lcout(N_347_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g2_1_0_LC_7_3_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g2_1_0_LC_7_3_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g2_1_0_LC_7_3_7.LUT_INIT=16'b0111011101110111;
    LogicCell40 un114_pixel_1_0_3__g2_1_0_LC_7_3_7 (
            .in0(N__15592),
            .in1(N__16024),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un114_pixel_1_0_3__g2_1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJPPPPD1_0_3_LC_7_4_0.C_ON=1'b0;
    defparam beamY_RNIJPPPPD1_0_3_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIJPPPPD1_0_3_LC_7_4_0.LUT_INIT=16'b0010010001000010;
    LogicCell40 beamY_RNIJPPPPD1_0_3_LC_7_4_0 (
            .in0(N__12264),
            .in1(N__12281),
            .in2(N__10686),
            .in3(N__10669),
            .lcout(),
            .ltout(font_un28_pixel_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_i_m2_LC_7_4_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_i_m2_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_i_m2_LC_7_4_1.LUT_INIT=16'b1110101100101000;
    LogicCell40 un114_pixel_1_0_3__g0_i_m2_LC_7_4_1 (
            .in0(N__10780),
            .in1(N__14954),
            .in2(N__10774),
            .in3(N__14269),
            .lcout(N_346_0_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_5_am_6_LC_7_4_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_5_am_6_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_5_am_6_LC_7_4_2.LUT_INIT=16'b1100011111111100;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_5_am_6_LC_7_4_2 (
            .in0(N__15591),
            .in1(N__15337),
            .in2(N__15816),
            .in3(N__16019),
            .lcout(),
            .ltout(un116_pixel_5_am_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_6_LC_7_4_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_6_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_6_LC_7_4_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_5_ns_6_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(N__14753),
            .in2(N__10771),
            .in3(N__11812),
            .lcout(N_379),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_0_LC_7_4_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_0_LC_7_4_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_0_LC_7_4_5.LUT_INIT=16'b0100000100101000;
    LogicCell40 un114_pixel_1_0_3__g0_0_LC_7_4_5 (
            .in0(N__12280),
            .in1(N__10768),
            .in2(N__10762),
            .in3(N__12263),
            .lcout(font_un28_pixel_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_1_2_LC_7_4_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_1_2_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_1_2_LC_7_4_6.LUT_INIT=16'b0111111101111100;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_2_ns_1_2_LC_7_4_6 (
            .in0(N__15590),
            .in1(N__15336),
            .in2(N__15815),
            .in3(N__16017),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un116_pixel_2_ns_1Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_2_LC_7_4_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_2_LC_7_4_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_2_LC_7_4_7.LUT_INIT=16'b1100000011100010;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_2_ns_2_LC_7_4_7 (
            .in0(N__16018),
            .in1(N__14752),
            .in2(N__10753),
            .in3(N__13418),
            .lcout(N_362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_1_2_LC_7_5_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_1_2_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_1_2_LC_7_5_0.LUT_INIT=16'b0001000111111111;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_5_ns_1_2_LC_7_5_0 (
            .in0(N__14741),
            .in1(N__15580),
            .in2(_gnd_net_),
            .in3(N__15334),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un116_pixel_5_ns_1Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_2_LC_7_5_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_2_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_2_LC_7_5_1.LUT_INIT=16'b1000001101000000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_5_ns_2_LC_7_5_1 (
            .in0(N__16021),
            .in1(N__14742),
            .in2(N__10750),
            .in3(N__15812),
            .lcout(un116_pixel_5_ns_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_5_ns_1_4_LC_7_5_2.C_ON=1'b0;
    defparam un116_pixel_5_ns_1_4_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam un116_pixel_5_ns_1_4_LC_7_5_2.LUT_INIT=16'b0011100000111100;
    LogicCell40 un116_pixel_5_ns_1_4_LC_7_5_2 (
            .in0(N__15586),
            .in1(N__15335),
            .in2(N__15817),
            .in3(N__16022),
            .lcout(),
            .ltout(un116_pixel_5_ns_1Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2L0T663_0_LC_7_5_3.C_ON=1'b0;
    defparam beamY_RNI2L0T663_0_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI2L0T663_0_LC_7_5_3.LUT_INIT=16'b0010000110101001;
    LogicCell40 beamY_RNI2L0T663_0_LC_7_5_3 (
            .in0(N__16023),
            .in1(N__14743),
            .in2(N__10840),
            .in3(N__13422),
            .lcout(beamY_RNI2L0T663Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIPU5VF83_1_LC_7_5_6.C_ON=1'b0;
    defparam beamY_RNIPU5VF83_1_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIPU5VF83_1_LC_7_5_6.LUT_INIT=16'b0000111101010011;
    LogicCell40 beamY_RNIPU5VF83_1_LC_7_5_6 (
            .in0(N__10837),
            .in1(N__10831),
            .in2(N__15012),
            .in3(N__13292),
            .lcout(),
            .ltout(un116_pixel_7_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIVU1O9R_1_LC_7_5_7.C_ON=1'b0;
    defparam beamY_RNIVU1O9R_1_LC_7_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIVU1O9R_1_LC_7_5_7.LUT_INIT=16'b1000111110000101;
    LogicCell40 beamY_RNIVU1O9R_1_LC_7_5_7 (
            .in0(N__13293),
            .in1(N__10786),
            .in2(N__10825),
            .in3(N__10822),
            .lcout(beamY_RNIVU1O9RZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI57H3N31_0_1_LC_7_6_0.C_ON=1'b0;
    defparam beamY_RNI57H3N31_0_1_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI57H3N31_0_1_LC_7_6_0.LUT_INIT=16'b1101000010000000;
    LogicCell40 beamY_RNI57H3N31_0_1_LC_7_6_0 (
            .in0(N__14901),
            .in1(N__11793),
            .in2(N__13306),
            .in3(N__10804),
            .lcout(),
            .ltout(beamY_RNI57H3N31_0Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1J75181_1_LC_7_6_1.C_ON=1'b0;
    defparam beamY_RNI1J75181_1_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI1J75181_1_LC_7_6_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 beamY_RNI1J75181_1_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(N__10816),
            .in2(N__10807),
            .in3(N__10795),
            .lcout(beamY_RNI1J75181Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI896FQ3_0_LC_7_6_2.C_ON=1'b0;
    defparam beamY_RNI896FQ3_0_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI896FQ3_0_LC_7_6_2.LUT_INIT=16'b0010111100100000;
    LogicCell40 beamY_RNI896FQ3_0_LC_7_6_2 (
            .in0(N__14217),
            .in1(N__11938),
            .in2(N__14759),
            .in3(N__11074),
            .lcout(beamY_RNI896FQ3Z0Z_0),
            .ltout(beamY_RNI896FQ3Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI57H3N31_1_LC_7_6_3.C_ON=1'b0;
    defparam beamY_RNI57H3N31_1_LC_7_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI57H3N31_1_LC_7_6_3.LUT_INIT=16'b1011100011111111;
    LogicCell40 beamY_RNI57H3N31_1_LC_7_6_3 (
            .in0(N__11794),
            .in1(N__14900),
            .in2(N__10798),
            .in3(N__13295),
            .lcout(beamY_RNI57H3N31Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIAK9BMC1_0_LC_7_6_4.C_ON=1'b0;
    defparam beamY_RNIAK9BMC1_0_LC_7_6_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIAK9BMC1_0_LC_7_6_4.LUT_INIT=16'b0001000110011001;
    LogicCell40 beamY_RNIAK9BMC1_0_LC_7_6_4 (
            .in0(N__15754),
            .in1(N__14630),
            .in2(_gnd_net_),
            .in3(N__15584),
            .lcout(),
            .ltout(un116_pixel_2_ns_1_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIGO5PPV_0_LC_7_6_5.C_ON=1'b0;
    defparam beamY_RNIGO5PPV_0_LC_7_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIGO5PPV_0_LC_7_6_5.LUT_INIT=16'b0000100000111010;
    LogicCell40 beamY_RNIGO5PPV_0_LC_7_6_5 (
            .in0(N__15296),
            .in1(N__15755),
            .in2(N__10789),
            .in3(N__13363),
            .lcout(beamY_RNIGO5PPVZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un114_pixel_3_i_m2_i_m2_6_LC_7_6_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un114_pixel_3_i_m2_i_m2_6_LC_7_6_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un114_pixel_3_i_m2_i_m2_6_LC_7_6_6.LUT_INIT=16'b1000110101100110;
    LogicCell40 un114_pixel_1_0_3__un114_pixel_3_i_m2_i_m2_6_LC_7_6_6 (
            .in0(N__15753),
            .in1(N__15295),
            .in2(N__14244),
            .in3(N__16020),
            .lcout(N_41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_7_6_7.C_ON=1'b0;
    defparam beamY_1_LC_7_6_7.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_7_6_7.LUT_INIT=16'b0100010001101100;
    LogicCell40 beamY_1_LC_7_6_7 (
            .in0(N__11026),
            .in1(N__14902),
            .in2(N__14702),
            .in3(N__10977),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11882),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_7_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_7_0 (
            .in0(_gnd_net_),
            .in1(N__13599),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_7_7_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_7_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__11139),
            .in2(N__10900),
            .in3(N__10912),
            .lcout(if_generate_plus_mult1_un68_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_7_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_7_2 (
            .in0(_gnd_net_),
            .in1(N__11125),
            .in2(N__15544),
            .in3(N__10909),
            .lcout(if_generate_plus_mult1_un68_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_7_7_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_7_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_7_7_3 (
            .in0(N__15249),
            .in1(N__11140),
            .in2(N__11116),
            .in3(N__10906),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_7_7_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_s_5_LC_7_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_s_5_LC_7_7_4 (
            .in0(_gnd_net_),
            .in1(N__11104),
            .in2(_gnd_net_),
            .in3(N__10903),
            .lcout(un5_rowlto2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_7_7_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_i_LC_7_7_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_i_LC_7_7_5 (
            .in0(N__11538),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_row_8_7_1_LC_7_7_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_row_8_7_1_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_row_8_7_1_LC_7_7_6.LUT_INIT=16'b0011001000110000;
    LogicCell40 un114_pixel_1_0_3__un4_row_8_7_1_LC_7_7_6 (
            .in0(N__15287),
            .in1(N__10890),
            .in2(N__15545),
            .in3(N__16016),
            .lcout(un114_pixel_1_0_3__un4_row_8_7Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_rowlto3_sbtinv_LC_7_7_7.C_ON=1'b0;
    defparam un5_rowlto3_sbtinv_LC_7_7_7.SEQ_MODE=4'b0000;
    defparam un5_rowlto3_sbtinv_LC_7_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_rowlto3_sbtinv_LC_7_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15492),
            .lcout(un5_rowlto3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__11537),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__11131),
            .in2(N__11092),
            .in3(N__11119),
            .lcout(if_generate_plus_mult1_un61_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(N__11353),
            .in2(N__12508),
            .in3(N__11107),
            .lcout(if_generate_plus_mult1_un61_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3 (
            .in0(N__15499),
            .in1(N__11091),
            .in2(N__11338),
            .in3(N__11098),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(N__11320),
            .in2(_gnd_net_),
            .in3(N__11095),
            .lcout(un5_rowlto3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_8_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12503),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__N_37_i_LC_7_9_0.C_ON=1'b1;
    defparam un114_pixel_1_0_3__N_37_i_LC_7_9_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__N_37_i_LC_7_9_0.LUT_INIT=16'b0001000100010001;
    LogicCell40 un114_pixel_1_0_3__N_37_i_LC_7_9_0 (
            .in0(N__15081),
            .in1(N__14030),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_37_i),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_9_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_9_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_9_1 (
            .in0(_gnd_net_),
            .in1(N__11290),
            .in2(N__11211),
            .in3(N__11077),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_9_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_9_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_9_2 (
            .in0(_gnd_net_),
            .in1(N__11257),
            .in2(N__11230),
            .in3(N__11251),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8BLE3_LC_7_9_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8BLE3_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8BLE3_LC_7_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8BLE3_LC_7_9_3 (
            .in0(N__11193),
            .in1(N__11248),
            .in2(N__11212),
            .in3(N__11242),
            .lcout(charx_if_generate_plus_mult1_un40_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un33_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_LC_7_9_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_LC_7_9_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_LC_7_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_LC_7_9_4 (
            .in0(_gnd_net_),
            .in1(N__11239),
            .in2(_gnd_net_),
            .in3(N__11233),
            .lcout(charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_9_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_9_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11225),
            .lcout(charx_if_generate_plus_mult1_un26_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_0_LC_7_9_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_0_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_0_LC_7_9_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_0_LC_7_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11192),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_10_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_10_0 (
            .in0(_gnd_net_),
            .in1(N__13858),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEB2_LC_7_10_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEB2_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEB2_LC_7_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEB2_LC_7_10_1 (
            .in0(_gnd_net_),
            .in1(N__11296),
            .in2(N__11157),
            .in3(N__11197),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEBZ0Z2),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLIT2_LC_7_10_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLIT2_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLIT2_LC_7_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLIT2_LC_7_10_2 (
            .in0(_gnd_net_),
            .in1(N__11194),
            .in2(N__11176),
            .in3(N__11167),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLITZ0Z2),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNIPCKK6_LC_7_10_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNIPCKK6_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNIPCKK6_LC_7_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNIPCKK6_LC_7_10_3 (
            .in0(N__11456),
            .in1(N__11164),
            .in2(N__11158),
            .in3(N__11143),
            .lcout(charx_if_generate_plus_mult1_un47_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_LC_7_10_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_LC_7_10_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_LC_7_10_4 (
            .in0(_gnd_net_),
            .in1(N__11305),
            .in2(_gnd_net_),
            .in3(N__11299),
            .lcout(charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_10_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_1_LC_7_10_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_1_LC_7_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14031),
            .lcout(charx_if_generate_plus_mult1_un33_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_7_10_6.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_7_10_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_0_LC_7_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_0_LC_7_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15065),
            .lcout(charx_if_generate_plus_mult1_un26_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_10_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_10_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_10_7.LUT_INIT=16'b0101010111111111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_10_7 (
            .in0(N__12896),
            .in1(N__14032),
            .in2(_gnd_net_),
            .in3(N__16153),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_11_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_11_0 (
            .in0(_gnd_net_),
            .in1(N__13868),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_11_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_11_1 (
            .in0(_gnd_net_),
            .in1(N__11284),
            .in2(N__11380),
            .in3(N__11278),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_2),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_11_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_11_2 (
            .in0(_gnd_net_),
            .in1(N__12832),
            .in2(N__11371),
            .in3(N__11275),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_3),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_11_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_11_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_11_3 (
            .in0(_gnd_net_),
            .in1(N__11272),
            .in2(N__11362),
            .in3(N__11263),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_4),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_0_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_0_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_11_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_11_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_11_4 (
            .in0(_gnd_net_),
            .in1(N__16152),
            .in2(_gnd_net_),
            .in3(N__11260),
            .lcout(column_1_if_generate_plus_mult1_un47_sum0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_7_11_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_2_LC_7_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_2_LC_7_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14038),
            .lcout(un5_visiblex_i_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_11_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_11_6.LUT_INIT=16'b1000100010001000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_11_6 (
            .in0(N__16138),
            .in1(N__12924),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(if_generate_plus_mult1_un47_sum_0_cry_3_ma),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_7_11_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_7_11_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_7_11_7.LUT_INIT=16'b0101010101100110;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_7_11_7 (
            .in0(N__16151),
            .in1(N__15077),
            .in2(N__12935),
            .in3(N__14039),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0 (
            .in0(_gnd_net_),
            .in1(N__11652),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1 (
            .in0(_gnd_net_),
            .in1(N__13033),
            .in2(N__12963),
            .in3(N__11341),
            .lcout(if_generate_plus_mult1_un54_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2 (
            .in0(_gnd_net_),
            .in1(N__13005),
            .in2(N__12991),
            .in3(N__11323),
            .lcout(if_generate_plus_mult1_un54_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3 (
            .in0(N__12499),
            .in1(N__11476),
            .in2(N__12964),
            .in3(N__11311),
            .lcout(column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4 (
            .in0(_gnd_net_),
            .in1(N__13018),
            .in2(_gnd_net_),
            .in3(N__11308),
            .lcout(if_generate_plus_mult1_un54_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_0_LC_7_12_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_0_LC_7_12_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_0_LC_7_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_0_LC_7_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11457),
            .lcout(charx_if_generate_plus_mult1_un40_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_12_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_12_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_12_6.LUT_INIT=16'b1001100111000011;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_12_6 (
            .in0(N__11485),
            .in1(N__13004),
            .in2(N__14134),
            .in3(N__16154),
            .lcout(),
            .ltout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_12_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_12_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_12_7.LUT_INIT=16'b0000111111110000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11479),
            .in3(N__12956),
            .lcout(if_generate_plus_mult1_un54_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_7_13_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_7_13_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_7_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_7_13_0 (
            .in0(_gnd_net_),
            .in1(N__11650),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0O3_LC_7_13_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0O3_LC_7_13_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0O3_LC_7_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0O3_LC_7_13_1 (
            .in0(_gnd_net_),
            .in1(N__11470),
            .in2(N__11412),
            .in3(N__11461),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0OZ0Z3),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCD16_LC_7_13_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCD16_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCD16_LC_7_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCD16_LC_7_13_2 (
            .in0(_gnd_net_),
            .in1(N__11458),
            .in2(N__11437),
            .in3(N__11425),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCDZ0Z16),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI8V4DD_LC_7_13_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI8V4DD_LC_7_13_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI8V4DD_LC_7_13_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI8V4DD_LC_7_13_3 (
            .in0(N__11604),
            .in1(N__11422),
            .in2(N__11413),
            .in3(N__11398),
            .lcout(charx_if_generate_plus_mult1_un54_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_LC_7_13_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_LC_7_13_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_LC_7_13_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_LC_7_13_4 (
            .in0(_gnd_net_),
            .in1(N__11395),
            .in2(_gnd_net_),
            .in3(N__11386),
            .lcout(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6),
            .ltout(charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_0_LC_7_13_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_0_LC_7_13_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_0_LC_7_13_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_0_LC_7_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11383),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_7_13_7.C_ON=1'b0;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_7_13_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_4_c_RNIP022_1_LC_7_13_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_4_c_RNIP022_1_LC_7_13_7 (
            .in0(N__11651),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0 (
            .in0(_gnd_net_),
            .in1(N__11545),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLM67_LC_7_14_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLM67_LC_7_14_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLM67_LC_7_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLM67_LC_7_14_1 (
            .in0(_gnd_net_),
            .in1(N__11614),
            .in2(N__11574),
            .in3(N__11608),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLMZ0Z67),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSA_LC_7_14_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSA_LC_7_14_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSA_LC_7_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSA_LC_7_14_2 (
            .in0(_gnd_net_),
            .in1(N__11605),
            .in2(N__11593),
            .in3(N__11584),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSAZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIGEUQ_LC_7_14_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIGEUQ_LC_7_14_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIGEUQ_LC_7_14_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIGEUQ_LC_7_14_3 (
            .in0(N__11700),
            .in1(N__11581),
            .in2(N__11575),
            .in3(N__11560),
            .lcout(charx_if_generate_plus_mult1_un61_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_LC_7_14_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_LC_7_14_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_LC_7_14_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_LC_7_14_4 (
            .in0(_gnd_net_),
            .in1(N__11557),
            .in2(_gnd_net_),
            .in3(N__11551),
            .lcout(charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_7_14_6.C_ON=1'b0;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_7_14_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_3_c_RNINT02_0_LC_7_14_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_3_c_RNINT02_0_LC_7_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11546),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_15_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_15_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_15_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_15_0 (
            .in0(_gnd_net_),
            .in1(N__13603),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRD_LC_7_15_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRD_LC_7_15_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRD_LC_7_15_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRD_LC_7_15_1 (
            .in0(_gnd_net_),
            .in1(N__11494),
            .in2(N__11682),
            .in3(N__11488),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRDZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0L_LC_7_15_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0L_LC_7_15_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0L_LC_7_15_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0L_LC_7_15_2 (
            .in0(_gnd_net_),
            .in1(N__11731),
            .in2(N__11701),
            .in3(N__11725),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0LZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGJ7MJ1_LC_7_15_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGJ7MJ1_LC_7_15_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGJ7MJ1_LC_7_15_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGJ7MJ1_LC_7_15_3 (
            .in0(N__13161),
            .in1(N__11722),
            .in2(N__11683),
            .in3(N__11716),
            .lcout(charx_if_generate_plus_mult1_un68_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_LC_7_15_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_LC_7_15_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_LC_7_15_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_LC_7_15_4 (
            .in0(_gnd_net_),
            .in1(N__11713),
            .in2(_gnd_net_),
            .in3(N__11707),
            .lcout(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0),
            .ltout(charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_0_LC_7_15_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_0_LC_7_15_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_0_LC_7_15_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_0_LC_7_15_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11704),
            .in3(_gnd_net_),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_0_LC_7_15_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_0_LC_7_15_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_0_LC_7_15_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_0_LC_7_15_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11696),
            .lcout(charx_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSyncZ0_LC_8_1_6.C_ON=1'b0;
    defparam VSyncZ0_LC_8_1_6.SEQ_MODE=4'b1000;
    defparam VSyncZ0_LC_8_1_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 VSyncZ0_LC_8_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12060),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11884),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_3_am_2_LC_8_3_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_3_am_2_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_3_am_2_LC_8_3_0.LUT_INIT=16'b1101000011100001;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_3_am_2_LC_8_3_0 (
            .in0(N__15808),
            .in1(N__15382),
            .in2(N__14776),
            .in3(N__16028),
            .lcout(un116_pixel_3_am_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_2_0_LC_8_4_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_2_0_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_2_0_LC_8_4_0.LUT_INIT=16'b0011000001101100;
    LogicCell40 un114_pixel_1_0_3__g0_2_0_LC_8_4_0 (
            .in0(N__13424),
            .in1(N__14757),
            .in2(N__15015),
            .in3(N__13228),
            .lcout(N_368_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_13_LC_8_4_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_13_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_13_LC_8_4_1.LUT_INIT=16'b1100000011001010;
    LogicCell40 un114_pixel_1_0_3__g0_13_LC_8_4_1 (
            .in0(N__16012),
            .in1(N__13045),
            .in2(N__14777),
            .in3(N__13423),
            .lcout(),
            .ltout(N_1556_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_11_LC_8_4_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_11_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_11_LC_8_4_2.LUT_INIT=16'b1101100011011000;
    LogicCell40 un114_pixel_1_0_3__g0_11_LC_8_4_2 (
            .in0(N__15003),
            .in1(N__14278),
            .in2(N__11782),
            .in3(_gnd_net_),
            .lcout(N_389_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_0_0_LC_8_4_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_0_0_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_0_0_LC_8_4_3.LUT_INIT=16'b0000111100110101;
    LogicCell40 un114_pixel_1_0_3__g0_0_0_LC_8_4_3 (
            .in0(N__11779),
            .in1(N__13213),
            .in2(N__11770),
            .in3(N__13303),
            .lcout(),
            .ltout(un114_pixel_1_0_3__font_un126_pixel_1_d_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_LC_8_4_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_LC_8_4_4.LUT_INIT=16'b1000111110000101;
    LogicCell40 un114_pixel_1_0_3__g0_LC_8_4_4 (
            .in0(N__13304),
            .in1(N__11761),
            .in2(N__11755),
            .in3(N__11752),
            .lcout(),
            .ltout(g0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_i_m2_0_LC_8_4_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_i_m2_0_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_i_m2_0_LC_8_4_5.LUT_INIT=16'b1111000011100100;
    LogicCell40 un114_pixel_1_0_3__g0_i_m2_0_LC_8_4_5 (
            .in0(N__14758),
            .in1(N__11746),
            .in2(N__11740),
            .in3(N__13305),
            .lcout(N_400),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__m18_0_m2_LC_8_4_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__m18_0_m2_LC_8_4_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__m18_0_m2_LC_8_4_6.LUT_INIT=16'b1011101101010101;
    LogicCell40 un114_pixel_1_0_3__m18_0_m2_LC_8_4_6 (
            .in0(N__15791),
            .in1(N__15589),
            .in2(_gnd_net_),
            .in3(N__15333),
            .lcout(N_36),
            .ltout(N_36_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_1_4_LC_8_4_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_1_4_LC_8_4_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_1_4_LC_8_4_7.LUT_INIT=16'b0000001011001110;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_1_4_LC_8_4_7 (
            .in0(N__16011),
            .in1(N__14751),
            .in2(N__11737),
            .in3(N__13234),
            .lcout(un116_pixel_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIC1MEAP2_1_LC_8_5_0.C_ON=1'b0;
    defparam beamY_RNIC1MEAP2_1_LC_8_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIC1MEAP2_1_LC_8_5_0.LUT_INIT=16'b1010111110100000;
    LogicCell40 beamY_RNIC1MEAP2_1_LC_8_5_0 (
            .in0(N__14461),
            .in1(_gnd_net_),
            .in2(N__13426),
            .in3(N__14800),
            .lcout(),
            .ltout(un116_pixel_3_ns_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNILBST4T2_1_LC_8_5_1.C_ON=1'b0;
    defparam beamY_RNILBST4T2_1_LC_8_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNILBST4T2_1_LC_8_5_1.LUT_INIT=16'b1000111110000101;
    LogicCell40 beamY_RNILBST4T2_1_LC_8_5_1 (
            .in0(N__14986),
            .in1(N__13432),
            .in2(N__11734),
            .in3(N__11806),
            .lcout(beamY_RNILBST4T2Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__N_315_i_i_a3_0_LC_8_5_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__N_315_i_i_a3_0_LC_8_5_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__N_315_i_i_a3_0_LC_8_5_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 un114_pixel_1_0_3__N_315_i_i_a3_0_LC_8_5_2 (
            .in0(_gnd_net_),
            .in1(N__15577),
            .in2(_gnd_net_),
            .in3(N__15326),
            .lcout(N_563),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_LC_8_5_3.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_LC_8_5_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_LC_8_5_3.LUT_INIT=16'b1010010111110000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_LC_8_5_3 (
            .in0(N__13543),
            .in1(_gnd_net_),
            .in2(N__13513),
            .in3(N__13464),
            .lcout(font_un3_pixel_29),
            .ltout(font_un3_pixel_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_7_x1_0_LC_8_5_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_7_x1_0_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_7_x1_0_LC_8_5_4.LUT_INIT=16'b0111111101001111;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_7_x1_0_LC_8_5_4 (
            .in0(N__13318),
            .in1(N__14987),
            .in2(N__11815),
            .in3(N__13334),
            .lcout(un116_pixel_7_x1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_5_bm_6_LC_8_5_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_5_bm_6_LC_8_5_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_5_bm_6_LC_8_5_5.LUT_INIT=16'b1001110010111110;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_5_bm_6_LC_8_5_5 (
            .in0(N__16000),
            .in1(N__15807),
            .in2(N__15384),
            .in3(N__14238),
            .lcout(un116_pixel_5_bm_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__m5_LC_8_5_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__m5_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__m5_LC_8_5_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 un114_pixel_1_0_3__m5_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(N__15578),
            .in2(_gnd_net_),
            .in3(N__15998),
            .lcout(N_325),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_4_bm_1_LC_8_5_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_4_bm_1_LC_8_5_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_4_bm_1_LC_8_5_7.LUT_INIT=16'b1101011011110110;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_4_bm_1_LC_8_5_7 (
            .in0(N__15999),
            .in1(N__15806),
            .in2(N__15383),
            .in3(N__15579),
            .lcout(un116_pixel_4_bm_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1C50FS3_0_LC_8_6_0.C_ON=1'b0;
    defparam beamY_RNI1C50FS3_0_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI1C50FS3_0_LC_8_6_0.LUT_INIT=16'b0000110011111010;
    LogicCell40 beamY_RNI1C50FS3_0_LC_8_6_0 (
            .in0(N__13381),
            .in1(N__13375),
            .in2(N__14775),
            .in3(N__14161),
            .lcout(),
            .ltout(beamY_RNI1C50FS3Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un126_pixel_2_bm_LC_8_6_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un126_pixel_2_bm_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un126_pixel_2_bm_LC_8_6_1.LUT_INIT=16'b1111000011001100;
    LogicCell40 un114_pixel_1_0_3__font_un126_pixel_2_bm_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(N__13204),
            .in2(N__11800),
            .in3(N__13300),
            .lcout(font_un126_pixel_2_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIG8FT9A2_0_LC_8_6_2.C_ON=1'b0;
    defparam beamY_RNIG8FT9A2_0_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIG8FT9A2_0_LC_8_6_2.LUT_INIT=16'b0100011100000101;
    LogicCell40 beamY_RNIG8FT9A2_0_LC_8_6_2 (
            .in0(N__15770),
            .in1(N__15588),
            .in2(N__14774),
            .in3(N__15288),
            .lcout(),
            .ltout(un116_pixel_3_bm_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIOHI2NG_0_LC_8_6_3.C_ON=1'b0;
    defparam beamY_RNIOHI2NG_0_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIOHI2NG_0_LC_8_6_3.LUT_INIT=16'b0101111101110100;
    LogicCell40 beamY_RNIOHI2NG_0_LC_8_6_3 (
            .in0(N__16009),
            .in1(N__14736),
            .in2(N__11797),
            .in3(N__15294),
            .lcout(beamY_RNIOHI2NGZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_0_LC_8_6_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_0_LC_8_6_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_2_ns_0_LC_8_6_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_2_ns_0_LC_8_6_4 (
            .in0(N__14737),
            .in1(N__13624),
            .in2(_gnd_net_),
            .in3(N__15442),
            .lcout(),
            .ltout(N_364_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI57H3N31_1_1_LC_8_6_5.C_ON=1'b0;
    defparam beamY_RNI57H3N31_1_1_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI57H3N31_1_1_LC_8_6_5.LUT_INIT=16'b0101010100100111;
    LogicCell40 beamY_RNI57H3N31_1_1_LC_8_6_5 (
            .in0(N__14903),
            .in1(N__13369),
            .in2(N__11950),
            .in3(N__13299),
            .lcout(),
            .ltout(un116_pixel_7_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI7OE17C_0_LC_8_6_6.C_ON=1'b0;
    defparam beamY_RNI7OE17C_0_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI7OE17C_0_LC_8_6_6.LUT_INIT=16'b1000111110000101;
    LogicCell40 beamY_RNI7OE17C_0_LC_8_6_6 (
            .in0(N__13301),
            .in1(N__14545),
            .in2(N__11947),
            .in3(N__11944),
            .lcout(beamY_RNI7OE17CZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__column_0111_1_0_LC_8_6_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__column_0111_1_0_LC_8_6_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__column_0111_1_0_LC_8_6_7.LUT_INIT=16'b0000000001010101;
    LogicCell40 un114_pixel_1_0_3__column_0111_1_0_LC_8_6_7 (
            .in0(N__16010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15769),
            .lcout(column_0111_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un126_pixel_6_am_LC_8_7_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un126_pixel_6_am_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un126_pixel_6_am_LC_8_7_0.LUT_INIT=16'b1110110101001000;
    LogicCell40 un114_pixel_1_0_3__font_un126_pixel_6_am_LC_8_7_0 (
            .in0(N__13541),
            .in1(N__13240),
            .in2(N__13465),
            .in3(N__11932),
            .lcout(),
            .ltout(font_un126_pixel_6_am_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_1_1_LC_8_7_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_1_1_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_1_1_LC_8_7_1.LUT_INIT=16'b0111001101100010;
    LogicCell40 un114_pixel_1_0_3__g0_1_1_LC_8_7_1 (
            .in0(N__12023),
            .in1(N__11821),
            .in2(N__11926),
            .in3(N__12127),
            .lcout(),
            .ltout(N_1075_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_4_LC_8_7_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_4_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_4_LC_8_7_2.LUT_INIT=16'b0101010001000100;
    LogicCell40 un114_pixel_1_0_3__g0_4_LC_8_7_2 (
            .in0(N__11923),
            .in1(N__12310),
            .in2(N__11911),
            .in3(N__12067),
            .lcout(),
            .ltout(Pixel_r_rn_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PixelZ0_LC_8_7_3.C_ON=1'b0;
    defparam PixelZ0_LC_8_7_3.SEQ_MODE=4'b1000;
    defparam PixelZ0_LC_8_7_3.LUT_INIT=16'b1100110011110000;
    LogicCell40 PixelZ0_LC_8_7_3 (
            .in0(_gnd_net_),
            .in1(N__11908),
            .in2(N__11899),
            .in3(N__12031),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__11883),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_7_LC_8_7_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_7_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_7_LC_8_7_4.LUT_INIT=16'b0010010101110101;
    LogicCell40 un114_pixel_1_0_3__g0_7_LC_8_7_4 (
            .in0(N__11839),
            .in1(N__11827),
            .in2(N__12025),
            .in3(N__13186),
            .lcout(un114_pixel_1_0_3__font_un126_pixel_7_d_ns_1_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI90K6F01_2_LC_8_7_5.C_ON=1'b0;
    defparam beamY_RNI90K6F01_2_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI90K6F01_2_LC_8_7_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 beamY_RNI90K6F01_2_LC_8_7_5 (
            .in0(_gnd_net_),
            .in1(N__12292),
            .in2(_gnd_net_),
            .in3(N__12265),
            .lcout(chary_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un126_pixel_6_bm_LC_8_7_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un126_pixel_6_bm_LC_8_7_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un126_pixel_6_bm_LC_8_7_6.LUT_INIT=16'b1111100101100000;
    LogicCell40 un114_pixel_1_0_3__font_un126_pixel_6_bm_LC_8_7_6 (
            .in0(N__13540),
            .in1(N__13460),
            .in2(N__12145),
            .in3(N__12136),
            .lcout(font_un126_pixel_6_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAV9A43_LC_8_8_0.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAV9A43_LC_8_8_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAV9A43_LC_8_8_0.LUT_INIT=16'b1100110000110011;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAV9A43_LC_8_8_0 (
            .in0(_gnd_net_),
            .in1(N__14451),
            .in2(_gnd_net_),
            .in3(N__13663),
            .lcout(charx_if_generate_plus_mult1_un1_sum_axb1),
            .ltout(charx_if_generate_plus_mult1_un1_sum_axb1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_0_LC_8_8_1.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_0_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_0_LC_8_8_1.LUT_INIT=16'b0000110000110000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_0_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__13509),
            .in2(N__12121),
            .in3(N__13458),
            .lcout(),
            .ltout(r_i1_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un126_pixel_m_2_LC_8_8_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un126_pixel_m_2_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un126_pixel_m_2_LC_8_8_2.LUT_INIT=16'b1000110001001100;
    LogicCell40 un114_pixel_1_0_3__font_un126_pixel_m_2_LC_8_8_2 (
            .in0(N__13492),
            .in1(N__12117),
            .in2(N__12094),
            .in3(N__12018),
            .lcout(),
            .ltout(un114_pixel_1_0_3__font_un126_pixel_mZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un126_pixel_m_1_LC_8_8_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un126_pixel_m_1_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un126_pixel_m_1_LC_8_8_3.LUT_INIT=16'b0110000000000000;
    LogicCell40 un114_pixel_1_0_3__font_un126_pixel_m_1_LC_8_8_3 (
            .in0(N__12360),
            .in1(N__12342),
            .in2(N__12091),
            .in3(N__12370),
            .lcout(),
            .ltout(un114_pixel_1_0_3__font_un126_pixel_m_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un126_pixel_m_3_LC_8_8_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un126_pixel_m_3_LC_8_8_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un126_pixel_m_3_LC_8_8_4.LUT_INIT=16'b1011000001100000;
    LogicCell40 un114_pixel_1_0_3__font_un126_pixel_m_3_LC_8_8_4 (
            .in0(N__14974),
            .in1(N__12088),
            .in2(N__12076),
            .in3(N__12073),
            .lcout(un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3),
            .ltout(un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_0_LC_8_8_5.C_ON=1'b0;
    defparam Pixel_RNO_0_LC_8_8_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_0_LC_8_8_5.LUT_INIT=16'b0001000000000000;
    LogicCell40 Pixel_RNO_0_LC_8_8_5 (
            .in0(N__12061),
            .in1(N__12306),
            .in2(N__12034),
            .in3(N__12826),
            .lcout(Pixel_r_sn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un57_pixel_0_LC_8_8_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un57_pixel_0_LC_8_8_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un57_pixel_0_LC_8_8_6.LUT_INIT=16'b0110011000000000;
    LogicCell40 un114_pixel_1_0_3__font_un57_pixel_0_LC_8_8_6 (
            .in0(N__13459),
            .in1(N__13542),
            .in2(_gnd_net_),
            .in3(N__12019),
            .lcout(un114_pixel_1_0_3__font_un57_pixelZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_row_8_3_LC_8_9_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_row_8_3_LC_8_9_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_row_8_3_LC_8_9_0.LUT_INIT=16'b1011000001010000;
    LogicCell40 un114_pixel_1_0_3__un4_row_8_3_LC_8_9_0 (
            .in0(N__12601),
            .in1(N__12820),
            .in2(N__12478),
            .in3(N__12691),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un4_row_8Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_row_8_7_LC_8_9_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_row_8_7_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_row_8_7_LC_8_9_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 un114_pixel_1_0_3__un4_row_8_7_LC_8_9_1 (
            .in0(N__12730),
            .in1(N__12447),
            .in2(N__12703),
            .in3(N__12700),
            .lcout(un114_pixel_1_0_3__un4_row_8Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_row_8_2_LC_8_9_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_row_8_2_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_row_8_2_LC_8_9_3.LUT_INIT=16'b0111000000000000;
    LogicCell40 un114_pixel_1_0_3__un4_row_8_2_LC_8_9_3 (
            .in0(N__12690),
            .in1(N__12600),
            .in2(N__12853),
            .in3(N__12507),
            .lcout(un114_pixel_1_0_3__un4_row_8Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_row_8_LC_8_9_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_row_8_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_row_8_LC_8_9_5.LUT_INIT=16'b0110100100000000;
    LogicCell40 un114_pixel_1_0_3__un4_row_8_LC_8_9_5 (
            .in0(N__12469),
            .in1(N__12448),
            .in2(N__12418),
            .in3(N__12376),
            .lcout(un114_pixel_1_0_3__un4_rowZ0Z_8),
            .ltout(un114_pixel_1_0_3__un4_rowZ0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__Pixel_3_sqmuxa_LC_8_9_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__Pixel_3_sqmuxa_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__Pixel_3_sqmuxa_LC_8_9_6.LUT_INIT=16'b1001111100000000;
    LogicCell40 un114_pixel_1_0_3__Pixel_3_sqmuxa_LC_8_9_6 (
            .in0(N__12364),
            .in1(N__12343),
            .in2(N__12322),
            .in3(N__12319),
            .lcout(Pixel_3_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_1_LC_8_9_7.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_1_LC_8_9_7.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_1_LC_8_9_7.LUT_INIT=16'b0100101111110000;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_1_LC_8_9_7 (
            .in0(N__14450),
            .in1(N__13719),
            .in2(N__13690),
            .in3(N__13659),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_10_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_10_0 (
            .in0(_gnd_net_),
            .in1(N__14425),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46K1_LC_8_10_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46K1_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46K1_LC_8_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46K1_LC_8_10_1 (
            .in0(_gnd_net_),
            .in1(N__12859),
            .in2(N__12841),
            .in3(N__12295),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9F2_LC_8_10_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9F2_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9F2_LC_8_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9F2_LC_8_10_2 (
            .in0(_gnd_net_),
            .in1(N__13177),
            .in2(N__13081),
            .in3(N__12877),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3 (
            .in0(_gnd_net_),
            .in1(N__13141),
            .in2(N__12874),
            .in3(N__13077),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_4_c_invZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPAC843_LC_8_10_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPAC843_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPAC843_LC_8_10_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPAC843_LC_8_10_4 (
            .in0(_gnd_net_),
            .in1(N__13105),
            .in2(_gnd_net_),
            .in3(N__12865),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843),
            .ltout(charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_8_10_5.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_8_10_5.LUT_INIT=16'b1010111101010000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_8_10_5 (
            .in0(N__14426),
            .in1(_gnd_net_),
            .in2(N__12862),
            .in3(N__13713),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_10_7.C_ON=1'b0;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15148),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_N_858_i_LC_8_11_0.C_ON=1'b0;
    defparam column_1_N_858_i_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam column_1_N_858_i_LC_8_11_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_N_858_i_LC_8_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16184),
            .lcout(N_858_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un4_row_8_0_LC_8_11_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un4_row_8_0_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un4_row_8_0_LC_8_11_1.LUT_INIT=16'b1101100001010000;
    LogicCell40 un114_pixel_1_0_3__un4_row_8_0_LC_8_11_1 (
            .in0(N__16186),
            .in1(N__12923),
            .in2(N__14098),
            .in3(N__12982),
            .lcout(un114_pixel_1_0_3__un4_row_8Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_0_LC_8_11_3.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_0_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_0_LC_8_11_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_0_LC_8_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13076),
            .lcout(charx_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_11_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_11_4.LUT_INIT=16'b1100011011111010;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_11_4 (
            .in0(N__14004),
            .in1(N__12919),
            .in2(N__12934),
            .in3(N__16185),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_6.LUT_INIT=16'b0001000111101110;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_6 (
            .in0(N__14003),
            .in1(N__12918),
            .in2(_gnd_net_),
            .in3(N__16183),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_sx_LC_8_12_0.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_sx_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_sx_LC_8_12_0.LUT_INIT=16'b0000100100001001;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_2_sx_LC_8_12_0 (
            .in0(N__13886),
            .in1(N__14089),
            .in2(N__16209),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(column_1_if_generate_plus_mult1_un54_sum_axb_2_sxZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_8_12_1.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_8_12_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_8_12_1.LUT_INIT=16'b0000011100001101;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_8_12_1 (
            .in0(N__16201),
            .in1(N__13887),
            .in2(N__13039),
            .in3(N__12981),
            .lcout(),
            .ltout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_8_12_2.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_8_12_2.LUT_INIT=16'b0000111111110000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_8_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13036),
            .in3(N__12955),
            .lcout(if_generate_plus_mult1_un54_sum_axb_2_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_8_12_3.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_m_5_LC_8_12_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_m_5_LC_8_12_3 (
            .in0(_gnd_net_),
            .in1(N__16191),
            .in2(N__14097),
            .in3(N__12979),
            .lcout(if_generate_plus_mult1_un47_sum_m_5),
            .ltout(if_generate_plus_mult1_un47_sum_m_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_8_12_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_8_12_4.LUT_INIT=16'b1100001110100101;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_8_12_4 (
            .in0(N__14110),
            .in1(N__13027),
            .in2(N__13021),
            .in3(N__16203),
            .lcout(column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_8_12_5.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_8_12_5.LUT_INIT=16'b1101100011011000;
    LogicCell40 column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_8_12_5 (
            .in0(N__16202),
            .in1(N__13012),
            .in2(N__13819),
            .in3(N__13006),
            .lcout(if_generate_plus_mult1_un54_sum_axb_3_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_N_584_i_LC_8_12_6.C_ON=1'b0;
    defparam column_1_N_584_i_LC_8_12_6.SEQ_MODE=4'b0000;
    defparam column_1_N_584_i_LC_8_12_6.LUT_INIT=16'b0101001101010011;
    LogicCell40 column_1_N_584_i_LC_8_12_6 (
            .in0(N__12980),
            .in1(N__14093),
            .in2(N__16208),
            .in3(_gnd_net_),
            .lcout(N_584_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_12_7.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_12_7.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_12_7.LUT_INIT=16'b0000110000111111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_12_7 (
            .in0(_gnd_net_),
            .in1(N__16190),
            .in2(N__14005),
            .in3(N__12936),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_14_0.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_14_0.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_14_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_14_0 (
            .in0(_gnd_net_),
            .in1(N__15155),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5R_LC_8_14_1.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5R_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5R_LC_8_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5R_LC_8_14_1 (
            .in0(_gnd_net_),
            .in1(N__13051),
            .in2(N__13119),
            .in3(N__13165),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5RZ0),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BV81_LC_8_14_2.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BV81_LC_8_14_2.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BV81_LC_8_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BV81_LC_8_14_2 (
            .in0(_gnd_net_),
            .in1(N__13162),
            .in2(N__13150),
            .in3(N__13129),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BVZ0Z81),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI3P7U33_LC_8_14_3.C_ON=1'b1;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI3P7U33_LC_8_14_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI3P7U33_LC_8_14_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI3P7U33_LC_8_14_3 (
            .in0(N__13070),
            .in1(N__13126),
            .in2(N__13120),
            .in3(N__13093),
            .lcout(charx_if_generate_plus_mult1_un75_sum_axb_5),
            .ltout(),
            .carryin(charx_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(charx_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_LC_8_14_4.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_LC_8_14_4.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_LC_8_14_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_LC_8_14_4 (
            .in0(_gnd_net_),
            .in1(N__13090),
            .in2(_gnd_net_),
            .in3(N__13084),
            .lcout(charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_8_14_7.C_ON=1'b0;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_8_14_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_2_c_RNILQV1_0_LC_8_14_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_2_c_RNILQV1_0_LC_8_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13611),
            .lcout(charx_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_i_m2_1_LC_9_4_0.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_i_m2_1_LC_9_4_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_i_m2_1_LC_9_4_0.LUT_INIT=16'b1010010101110010;
    LogicCell40 un114_pixel_1_0_3__g0_i_m2_1_LC_9_4_0 (
            .in0(N__16002),
            .in1(N__14239),
            .in2(N__15405),
            .in3(N__15793),
            .lcout(N_41_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g1_4_LC_9_4_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g1_4_LC_9_4_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g1_4_LC_9_4_1.LUT_INIT=16'b1010101001010101;
    LogicCell40 un114_pixel_1_0_3__g1_4_LC_9_4_1 (
            .in0(N__15795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15608),
            .lcout(un114_pixel_1_0_3__g1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__column_0111_0_LC_9_4_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__column_0111_0_LC_9_4_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__column_0111_0_LC_9_4_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 un114_pixel_1_0_3__column_0111_0_LC_9_4_3 (
            .in0(N__15792),
            .in1(N__15385),
            .in2(_gnd_net_),
            .in3(N__16001),
            .lcout(column_0111_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_3_1_LC_9_4_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_3_1_LC_9_4_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_3_1_LC_9_4_5.LUT_INIT=16'b0000001011110001;
    LogicCell40 un114_pixel_1_0_3__g0_3_1_LC_9_4_5 (
            .in0(N__15796),
            .in1(N__15389),
            .in2(N__15014),
            .in3(N__16003),
            .lcout(un116_pixel_3_ns_1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_17_LC_9_4_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_17_LC_9_4_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_17_LC_9_4_6.LUT_INIT=16'b1010111101110010;
    LogicCell40 un114_pixel_1_0_3__g0_17_LC_9_4_6 (
            .in0(N__16004),
            .in1(N__14240),
            .in2(N__15406),
            .in3(N__15794),
            .lcout(),
            .ltout(N_1583_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_14_LC_9_4_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_14_LC_9_4_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_14_LC_9_4_7.LUT_INIT=16'b1110010010100000;
    LogicCell40 un114_pixel_1_0_3__g0_14_LC_9_4_7 (
            .in0(N__14999),
            .in1(N__13222),
            .in2(N__13216),
            .in3(N__15393),
            .lcout(N_26_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_2_am_1_LC_9_5_0.C_ON=1'b0;
    defparam un116_pixel_2_am_1_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam un116_pixel_2_am_1_LC_9_5_0.LUT_INIT=16'b1000101101000100;
    LogicCell40 un116_pixel_2_am_1_LC_9_5_0 (
            .in0(N__15395),
            .in1(N__15804),
            .in2(N__14254),
            .in3(N__16007),
            .lcout(),
            .ltout(un116_pixel_2_amZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_6_1_LC_9_5_1.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_6_1_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_6_1_LC_9_5_1.LUT_INIT=16'b1101100111001000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_6_1_LC_9_5_1 (
            .in0(N__14985),
            .in1(N__13345),
            .in2(N__13207),
            .in3(N__13351),
            .lcout(un116_pixel_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_4_0_15__m15_0_a3_LC_9_5_2.C_ON=1'b0;
    defparam un114_pixel_4_0_15__m15_0_a3_LC_9_5_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_4_0_15__m15_0_a3_LC_9_5_2.LUT_INIT=16'b0010001000000000;
    LogicCell40 un114_pixel_4_0_15__m15_0_a3_LC_9_5_2 (
            .in0(N__14237),
            .in1(N__15805),
            .in2(_gnd_net_),
            .in3(N__16008),
            .lcout(),
            .ltout(column_0001_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIT81CMJ2_1_LC_9_5_3.C_ON=1'b0;
    defparam beamY_RNIT81CMJ2_1_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIT81CMJ2_1_LC_9_5_3.LUT_INIT=16'b1111011110100010;
    LogicCell40 beamY_RNIT81CMJ2_1_LC_9_5_3 (
            .in0(N__14984),
            .in1(N__14746),
            .in2(N__13198),
            .in3(N__13335),
            .lcout(),
            .ltout(beamY_RNIT81CMJ2Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__font_un126_pixel_2_am_LC_9_5_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__font_un126_pixel_2_am_LC_9_5_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__font_un126_pixel_2_am_LC_9_5_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 un114_pixel_1_0_3__font_un126_pixel_2_am_LC_9_5_4 (
            .in0(_gnd_net_),
            .in1(N__13195),
            .in2(N__13189),
            .in3(N__13294),
            .lcout(font_un126_pixel_2_am),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_4_am_1_LC_9_5_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_4_am_1_LC_9_5_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_4_am_1_LC_9_5_6.LUT_INIT=16'b1101000110111011;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_4_am_1_LC_9_5_6 (
            .in0(N__15394),
            .in1(N__15803),
            .in2(N__14253),
            .in3(N__16005),
            .lcout(un116_pixel_4_am_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__m20_LC_9_5_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__m20_LC_9_5_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__m20_LC_9_5_7.LUT_INIT=16'b1100110001000100;
    LogicCell40 un114_pixel_1_0_3__m20_LC_9_5_7 (
            .in0(N__16006),
            .in1(N__14745),
            .in2(_gnd_net_),
            .in3(N__13425),
            .lcout(N_374_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_5_am_5_LC_9_6_0.C_ON=1'b0;
    defparam un116_pixel_5_am_5_LC_9_6_0.SEQ_MODE=4'b0000;
    defparam un116_pixel_5_am_5_LC_9_6_0.LUT_INIT=16'b0101101010001000;
    LogicCell40 un116_pixel_5_am_5_LC_9_6_0 (
            .in0(N__16014),
            .in1(N__14221),
            .in2(N__15404),
            .in3(N__15757),
            .lcout(un116_pixel_5_amZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_2_am_5_LC_9_6_1.C_ON=1'b0;
    defparam un116_pixel_2_am_5_LC_9_6_1.SEQ_MODE=4'b0000;
    defparam un116_pixel_2_am_5_LC_9_6_1.LUT_INIT=16'b1100000011010001;
    LogicCell40 un116_pixel_2_am_5_LC_9_6_1 (
            .in0(N__15758),
            .in1(N__16015),
            .in2(N__14246),
            .in3(N__15380),
            .lcout(un116_pixel_2_amZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_0_LC_9_6_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_0_LC_9_6_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_0_LC_9_6_2.LUT_INIT=16'b1111011111000000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_5_ns_0_LC_9_6_2 (
            .in0(N__15381),
            .in1(N__13618),
            .in2(N__14773),
            .in3(N__15760),
            .lcout(N_385),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_2_bm_1_LC_9_6_3.C_ON=1'b0;
    defparam un116_pixel_2_bm_1_LC_9_6_3.SEQ_MODE=4'b0000;
    defparam un116_pixel_2_bm_1_LC_9_6_3.LUT_INIT=16'b1100110011101110;
    LogicCell40 un116_pixel_2_bm_1_LC_9_6_3 (
            .in0(N__15759),
            .in1(N__13362),
            .in2(_gnd_net_),
            .in3(N__15375),
            .lcout(un116_pixel_2_bmZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_6_1_1_LC_9_6_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_6_1_1_LC_9_6_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_6_1_1_LC_9_6_4.LUT_INIT=16'b1111010110000101;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_6_1_1_LC_9_6_4 (
            .in0(N__14729),
            .in1(N__13552),
            .in2(N__14975),
            .in3(N__15761),
            .lcout(un114_pixel_1_0_3__un116_pixel_6_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_7_x0_0_LC_9_6_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_7_x0_0_LC_9_6_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_7_x0_0_LC_9_6_5.LUT_INIT=16'b0011101000000000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_7_x0_0_LC_9_6_5 (
            .in0(N__13339),
            .in1(N__13317),
            .in2(N__14976),
            .in3(N__13302),
            .lcout(),
            .ltout(un116_pixel_7_x0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_7_ns_0_LC_9_6_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_7_ns_0_LC_9_6_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_7_ns_0_LC_9_6_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_7_ns_0_LC_9_6_6 (
            .in0(_gnd_net_),
            .in1(N__14473),
            .in2(N__13249),
            .in3(N__13246),
            .lcout(un116_pixel_7_ns_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_2_bm_0_LC_9_6_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_2_bm_0_LC_9_6_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_2_bm_0_LC_9_6_7.LUT_INIT=16'b1000000011100110;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_2_bm_0_LC_9_6_7 (
            .in0(N__15756),
            .in1(N__16013),
            .in2(N__14245),
            .in3(N__15376),
            .lcout(un116_pixel_2_bm_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_1_0_0_LC_9_7_3.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_1_0_0_LC_9_7_3.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_5_ns_1_0_0_LC_9_7_3.LUT_INIT=16'b0101001111010011;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_5_ns_1_0_0_LC_9_7_3 (
            .in0(N__15594),
            .in1(N__15919),
            .in2(N__14744),
            .in3(N__15302),
            .lcout(un114_pixel_1_0_3__un116_pixel_5_ns_1_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_9_7_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un68_sum_i_LC_9_7_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un68_sum_i_LC_9_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13607),
            .lcout(column_1_if_generate_plus_mult1_un68_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_6_1_1_1_LC_9_7_7.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_6_1_1_1_LC_9_7_7.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_6_1_1_1_LC_9_7_7.LUT_INIT=16'b0101010111011101;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_6_1_1_1_LC_9_7_7 (
            .in0(N__15593),
            .in1(N__15918),
            .in2(_gnd_net_),
            .in3(N__15301),
            .lcout(un114_pixel_1_0_3__un116_pixel_6_1_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_8_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_8_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_8_0 (
            .in0(_gnd_net_),
            .in1(N__13536),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSO4_LC_9_8_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSO4_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSO4_LC_9_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSO4_LC_9_8_1 (
            .in0(_gnd_net_),
            .in1(N__13749),
            .in2(N__13729),
            .in3(N__13495),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3E987_LC_9_8_2.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3E987_LC_9_8_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3E987_LC_9_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3E987_LC_9_8_2 (
            .in0(_gnd_net_),
            .in1(N__13798),
            .in2(N__13482),
            .in3(N__13486),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3EZ0Z987),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_8_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_8_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_8_3 (
            .in0(_gnd_net_),
            .in1(N__13750),
            .in2(N__13789),
            .in3(N__13748),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CI987_LC_9_8_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CI987_LC_9_8_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CI987_LC_9_8_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CI987_LC_9_8_4 (
            .in0(N__13776),
            .in1(N__13762),
            .in2(N__13483),
            .in3(N__13468),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13807),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8T77_LC_9_9_1.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8T77_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8T77_LC_9_9_1.LUT_INIT=16'b1010010101011010;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8T77_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13633),
            .in3(N__13792),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8TZ0Z77),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(N__16397),
            .in2(N__13738),
            .in3(N__13780),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3.C_ON=1'b1;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13777),
            .in3(N__13756),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO),
            .ltout(),
            .carryin(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3),
            .carryout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4.C_ON=1'b0;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13753),
            .lcout(font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_0_LC_9_9_5.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_0_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_0_LC_9_9_5.LUT_INIT=16'b1011010000001111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_0_LC_9_9_5 (
            .in0(N__14445),
            .in1(N__13715),
            .in2(N__13689),
            .in3(N__13657),
            .lcout(charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIOUEGO4_LC_9_9_6.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIOUEGO4_LC_9_9_6.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIOUEGO4_LC_9_9_6.LUT_INIT=16'b0000111110100101;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIOUEGO4_LC_9_9_6 (
            .in0(N__13658),
            .in1(_gnd_net_),
            .in2(N__13720),
            .in3(N__14446),
            .lcout(charx_i_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_LC_9_10_3.C_ON=1'b0;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_LC_9_10_3.LUT_INIT=16'b1011010000001111;
    LogicCell40 charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_LC_9_10_3 (
            .in0(N__14444),
            .in1(N__13714),
            .in2(N__13688),
            .in3(N__13656),
            .lcout(charx_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_11_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(N__13888),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUH2_LC_9_11_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUH2_LC_9_11_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUH2_LC_9_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUH2_LC_9_11_1 (
            .in0(_gnd_net_),
            .in1(N__13894),
            .in2(N__14073),
            .in3(N__13948),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUHZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV6153_LC_9_11_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV6153_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV6153_LC_9_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV6153_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(N__14365),
            .in2(N__13984),
            .in3(N__13933),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIVZ0Z6153),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNISAMG7_LC_9_11_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNISAMG7_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNISAMG7_LC_9_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNISAMG7_LC_9_11_3 (
            .in0(N__13910),
            .in1(N__13969),
            .in2(N__14074),
            .in3(N__13921),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_LC_9_11_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_LC_9_11_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_LC_9_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_LC_9_11_4 (
            .in0(_gnd_net_),
            .in1(N__14380),
            .in2(_gnd_net_),
            .in3(N__13918),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_9_11_5.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_9_11_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_3_LC_9_11_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_3_LC_9_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14057),
            .lcout(un5_visiblex_i_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_9_11_7.C_ON=1'b0;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_9_11_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_6_c_RNIT642_0_LC_9_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_6_c_RNIT642_0_LC_9_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14058),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_9_12_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_9_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_9_12_0 (
            .in0(_gnd_net_),
            .in1(N__13885),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_9_12_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_9_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_9_12_1 (
            .in0(_gnd_net_),
            .in1(N__16198),
            .in2(N__13828),
            .in3(N__13810),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_2),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_9_12_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_9_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_9_12_2 (
            .in0(_gnd_net_),
            .in1(N__14149),
            .in2(N__14143),
            .in3(N__14122),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_3),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_9_12_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_9_12_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_9_12_3 (
            .in0(_gnd_net_),
            .in1(N__16199),
            .in2(N__14119),
            .in3(N__14104),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_4),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un47_sum_1_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un47_sum_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_9_12_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_9_12_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_9_12_4.LUT_INIT=16'b1000000001111111;
    LogicCell40 column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_9_12_4 (
            .in0(N__16200),
            .in1(N__14059),
            .in2(N__15106),
            .in3(N__14101),
            .lcout(column_1_if_generate_plus_mult1_un47_sum1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_0_LC_9_12_5.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_0_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_0_LC_9_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_0_LC_9_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14360),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_0_LC_9_12_6.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_0_LC_9_12_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_0_LC_9_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_0_LC_9_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16236),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__SUM4_3_i_a2_LC_9_13_0.C_ON=1'b1;
    defparam un114_pixel_1_0_3__SUM4_3_i_a2_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__SUM4_3_i_a2_LC_9_13_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 un114_pixel_1_0_3__SUM4_3_i_a2_LC_9_13_0 (
            .in0(_gnd_net_),
            .in1(N__14048),
            .in2(_gnd_net_),
            .in3(N__15097),
            .lcout(N_66),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5L_LC_9_13_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5L_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5L_LC_9_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5L_LC_9_13_1 (
            .in0(_gnd_net_),
            .in1(N__14388),
            .in2(N__14344),
            .in3(N__13972),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5LZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7J31_LC_9_13_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7J31_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7J31_LC_9_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7J31_LC_9_13_2 (
            .in0(_gnd_net_),
            .in1(N__16240),
            .in2(N__16429),
            .in3(N__13960),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7JZ0Z31),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8U9I3_LC_9_13_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8U9I3_LC_9_13_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8U9I3_LC_9_13_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8U9I3_LC_9_13_3 (
            .in0(N__14361),
            .in1(N__14389),
            .in2(N__16276),
            .in3(N__14371),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_LC_9_13_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_LC_9_13_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_LC_9_13_4 (
            .in0(_gnd_net_),
            .in1(N__16258),
            .in2(_gnd_net_),
            .in3(N__14368),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_9_13_7.C_ON=1'b0;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_7_c_RNIV952_1_LC_9_13_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_visiblex_cry_7_c_RNIV952_1_LC_9_13_7 (
            .in0(N__15098),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_11_1_4.C_ON=1'b0;
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_11_1_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_11_1_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_11_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14335),
            .lcout(GB_BUFFER_Clock12MHz_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_15_LC_11_4_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_15_LC_11_4_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_15_LC_11_4_2.LUT_INIT=16'b0100000000011001;
    LogicCell40 un114_pixel_1_0_3__g0_15_LC_11_4_2 (
            .in0(N__15402),
            .in1(N__15789),
            .in2(N__14779),
            .in3(N__15996),
            .lcout(N_1557_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIKBQK731_0_LC_11_4_3.C_ON=1'b0;
    defparam beamY_RNIKBQK731_0_LC_11_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIKBQK731_0_LC_11_4_3.LUT_INIT=16'b0001000111111111;
    LogicCell40 beamY_RNIKBQK731_0_LC_11_4_3 (
            .in0(N__14769),
            .in1(N__15616),
            .in2(_gnd_net_),
            .in3(N__15401),
            .lcout(un116_pixel_2_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__g0_i_m2_2_LC_11_4_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__g0_i_m2_2_LC_11_4_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__g0_i_m2_2_LC_11_4_6.LUT_INIT=16'b1000101101100110;
    LogicCell40 un114_pixel_1_0_3__g0_i_m2_2_LC_11_4_6 (
            .in0(N__15403),
            .in1(N__15790),
            .in2(N__14260),
            .in3(N__15997),
            .lcout(N_41_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_5_bm_5_LC_11_5_0.C_ON=1'b0;
    defparam un116_pixel_5_bm_5_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam un116_pixel_5_bm_5_LC_11_5_0.LUT_INIT=16'b0111010000000000;
    LogicCell40 un116_pixel_5_bm_5_LC_11_5_0 (
            .in0(N__15397),
            .in1(N__15693),
            .in2(N__14256),
            .in3(N__15982),
            .lcout(),
            .ltout(un116_pixel_5_bmZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJEPU0R2_1_LC_11_5_1.C_ON=1'b0;
    defparam beamY_RNIJEPU0R2_1_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIJEPU0R2_1_LC_11_5_1.LUT_INIT=16'b0001100101011101;
    LogicCell40 beamY_RNIJEPU0R2_1_LC_11_5_1 (
            .in0(N__15010),
            .in1(N__14766),
            .in2(N__14164),
            .in3(N__14491),
            .lcout(un116_pixel_6_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__m33_LC_11_5_2.C_ON=1'b0;
    defparam un114_pixel_1_0_3__m33_LC_11_5_2.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__m33_LC_11_5_2.LUT_INIT=16'b0110010000010001;
    LogicCell40 un114_pixel_1_0_3__m33_LC_11_5_2 (
            .in0(N__15398),
            .in1(N__15695),
            .in2(N__15618),
            .in3(N__15983),
            .lcout(un114_pixel_6_1_5__N_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_2_bm_5_LC_11_5_3.C_ON=1'b0;
    defparam un116_pixel_2_bm_5_LC_11_5_3.SEQ_MODE=4'b0000;
    defparam un116_pixel_2_bm_5_LC_11_5_3.LUT_INIT=16'b0111011111111111;
    LogicCell40 un116_pixel_2_bm_5_LC_11_5_3 (
            .in0(N__15692),
            .in1(N__15609),
            .in2(_gnd_net_),
            .in3(N__15396),
            .lcout(un116_pixel_2_bmZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__m24_LC_11_5_4.C_ON=1'b0;
    defparam un114_pixel_1_0_3__m24_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__m24_LC_11_5_4.LUT_INIT=16'b0010000010011001;
    LogicCell40 un114_pixel_1_0_3__m24_LC_11_5_4 (
            .in0(N__15399),
            .in1(N__15694),
            .in2(N__15619),
            .in3(N__15984),
            .lcout(),
            .ltout(un114_pixel_7_1_7__N_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_1_0_LC_11_5_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_1_0_LC_11_5_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_1_0_LC_11_5_5.LUT_INIT=16'b0000110000011101;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_3_ns_1_0_LC_11_5_5 (
            .in0(N__15696),
            .in1(N__14767),
            .in2(N__14485),
            .in3(N__15400),
            .lcout(),
            .ltout(un114_pixel_1_0_3__un116_pixel_3_ns_1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_0_LC_11_5_6.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_0_LC_11_5_6.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_3_ns_0_LC_11_5_6.LUT_INIT=16'b0100001011011011;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_3_ns_0_LC_11_5_6 (
            .in0(N__14768),
            .in1(N__15011),
            .in2(N__14482),
            .in3(N__14479),
            .lcout(N_371),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJUCG3J3_1_LC_11_5_7.C_ON=1'b0;
    defparam beamY_RNIJUCG3J3_1_LC_11_5_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIJUCG3J3_1_LC_11_5_7.LUT_INIT=16'b0010001001100110;
    LogicCell40 beamY_RNIJUCG3J3_1_LC_11_5_7 (
            .in0(N__15009),
            .in1(N__14765),
            .in2(_gnd_net_),
            .in3(N__15022),
            .lcout(beamY_RNIJUCG3J3Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_11_6_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_11_6_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_11_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_11_6_0 (
            .in0(_gnd_net_),
            .in1(N__14452),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_11_6_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_11_6_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_11_6_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_11_6_1 (
            .in0(_gnd_net_),
            .in1(N__14395),
            .in2(N__15121),
            .in3(N__15861),
            .lcout(G_345),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_11_6_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_11_6_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_11_6_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_11_6_2 (
            .in0(_gnd_net_),
            .in1(N__14524),
            .in2(N__15917),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_11_6_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_11_6_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_11_6_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_11_6_3 (
            .in0(_gnd_net_),
            .in1(N__15034),
            .in2(N__14503),
            .in3(N__15862),
            .lcout(G_346),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un82_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un82_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_11_6_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_11_6_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_s_5_LC_11_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_s_5_LC_11_6_4 (
            .in0(_gnd_net_),
            .in1(N__16051),
            .in2(_gnd_net_),
            .in3(N__15028),
            .lcout(un5_rowlto0),
            .ltout(un5_rowlto0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un116_pixel_1_bm_1_LC_11_6_5.C_ON=1'b0;
    defparam un116_pixel_1_bm_1_LC_11_6_5.SEQ_MODE=4'b0000;
    defparam un116_pixel_1_bm_1_LC_11_6_5.LUT_INIT=16'b1000100011000011;
    LogicCell40 un116_pixel_1_bm_1_LC_11_6_5 (
            .in0(N__15587),
            .in1(N__15356),
            .in2(N__15025),
            .in3(N__15866),
            .lcout(un116_pixel_1_bmZ0Z_1),
            .ltout(un116_pixel_1_bmZ0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIV622TR_1_LC_11_6_6.C_ON=1'b0;
    defparam beamY_RNIV622TR_1_LC_11_6_6.SEQ_MODE=4'b0000;
    defparam beamY_RNIV622TR_1_LC_11_6_6.LUT_INIT=16'b0000001111101110;
    LogicCell40 beamY_RNIV622TR_1_LC_11_6_6 (
            .in0(N__15867),
            .in1(N__14920),
            .in2(N__14803),
            .in3(N__14761),
            .lcout(beamY_RNIV622TRZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIITCG3J3_0_LC_11_6_7.C_ON=1'b0;
    defparam beamY_RNIITCG3J3_0_LC_11_6_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIITCG3J3_0_LC_11_6_7.LUT_INIT=16'b0111000111010000;
    LogicCell40 beamY_RNIITCG3J3_0_LC_11_6_7 (
            .in0(N__15728),
            .in1(N__14788),
            .in2(N__14778),
            .in3(N__15868),
            .lcout(beamY_RNIITCG3J3Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_7_0.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_7_0.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_7_0 (
            .in0(_gnd_net_),
            .in1(N__15162),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_7_1.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_7_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_7_1 (
            .in0(_gnd_net_),
            .in1(N__15169),
            .in2(N__14536),
            .in3(N__14518),
            .lcout(if_generate_plus_mult1_un75_sum_cry_2_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_7_2.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_7_2.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_7_2 (
            .in0(_gnd_net_),
            .in1(N__15300),
            .in2(N__14515),
            .in3(N__14494),
            .lcout(if_generate_plus_mult1_un75_sum_cry_3_s),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_7_3.C_ON=1'b1;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_7_3.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_7_3 (
            .in0(N__15869),
            .in1(N__15412),
            .in2(N__15430),
            .in3(N__16045),
            .lcout(column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5),
            .ltout(),
            .carryin(column_1_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(column_1_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_7_4.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_7_4.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_7_4 (
            .in0(_gnd_net_),
            .in1(N__16042),
            .in2(_gnd_net_),
            .in3(N__16033),
            .lcout(un5_rowlto1),
            .ltout(un5_rowlto1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un114_pixel_1_0_3__un116_pixel_2_am_0_LC_11_7_5.C_ON=1'b0;
    defparam un114_pixel_1_0_3__un116_pixel_2_am_0_LC_11_7_5.SEQ_MODE=4'b0000;
    defparam un114_pixel_1_0_3__un116_pixel_2_am_0_LC_11_7_5.LUT_INIT=16'b1001111011011110;
    LogicCell40 un114_pixel_1_0_3__un116_pixel_2_am_0_LC_11_7_5 (
            .in0(N__15684),
            .in1(N__15299),
            .in2(N__15622),
            .in3(N__15617),
            .lcout(un116_pixel_2_am_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_7_6.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_7_6.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_7_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_7_6 (
            .in0(N__15298),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15429),
            .lcout(if_generate_plus_mult1_un75_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_rowlto2_sbtinv_LC_11_7_7.C_ON=1'b0;
    defparam un5_rowlto2_sbtinv_LC_11_7_7.SEQ_MODE=4'b0000;
    defparam un5_rowlto2_sbtinv_LC_11_7_7.LUT_INIT=16'b0011001100110011;
    LogicCell40 un5_rowlto2_sbtinv_LC_11_7_7 (
            .in0(_gnd_net_),
            .in1(N__15297),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_rowlto2_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_1.C_ON=1'b0;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_1.SEQ_MODE=4'b0000;
    defparam column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15163),
            .lcout(column_1_if_generate_plus_mult1_un75_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_11_11_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_11_11_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_11_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_11_11_0 (
            .in0(_gnd_net_),
            .in1(N__16207),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_11_1.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_11_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15109),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_12_0.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_12_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_12_0 (
            .in0(_gnd_net_),
            .in1(N__15102),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHG_LC_11_12_1.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHG_LC_11_12_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHG_LC_11_12_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHG_LC_11_12_1 (
            .in0(_gnd_net_),
            .in1(N__16081),
            .in2(_gnd_net_),
            .in3(N__16414),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHGZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6Q_LC_11_12_2.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6Q_LC_11_12_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6Q_LC_11_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6Q_LC_11_12_2 (
            .in0(_gnd_net_),
            .in1(N__16216),
            .in2(N__16411),
            .in3(N__16261),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6QZ0),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNITTA02_LC_11_12_3.C_ON=1'b1;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNITTA02_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNITTA02_LC_11_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNITTA02_LC_11_12_3 (
            .in0(N__16235),
            .in1(N__16075),
            .in2(N__16060),
            .in3(N__16246),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_LC_11_12_4.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_LC_11_12_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_LC_11_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_LC_11_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16243),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_11_12_5.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_11_12_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_11_12_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_11_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16072),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_11_12_6.C_ON=1'b0;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_11_12_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_cry_8_c_RNI1D62_0_LC_11_12_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_cry_8_c_RNI1D62_0_LC_11_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16210),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKN_LC_11_12_7.C_ON=1'b0;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKN_LC_11_12_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKN_LC_11_12_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKN_LC_11_12_7 (
            .in0(_gnd_net_),
            .in1(N__16073),
            .in2(_gnd_net_),
            .in3(N__16074),
            .lcout(chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKNZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
