-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 17 2015 18:20:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4260\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3492\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3453\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3231\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3213\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3147\ : std_logic;
signal \N__3144\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3120\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3063\ : std_logic;
signal \N__3060\ : std_logic;
signal \N__3057\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3042\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2997\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2887\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2871\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2854\ : std_logic;
signal \N__2851\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2793\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2681\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2675\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2664\ : std_logic;
signal \N__2661\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2643\ : std_logic;
signal \N__2634\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2606\ : std_logic;
signal \N__2603\ : std_logic;
signal \N__2600\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2568\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2562\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2556\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2522\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2477\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2465\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2442\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2388\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2342\ : std_logic;
signal \N__2339\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \VCCG0\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_7_1_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\ : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOMZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPMZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\ : std_logic;
signal \un5_visibley_cry_7_c_RNI1L4CZ0Z_0\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal \beamY_RNO_0Z0Z_3\ : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal \beamY_RNO_0Z0Z_4\ : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal \beamY_RNO_0Z0Z_7\ : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \beamY_RNO_0Z0Z_9\ : std_logic;
signal \un3_beamx_5_cascade_\ : std_logic;
signal un3_beamx_7 : std_logic;
signal \beamY_RNO_0Z0Z_1\ : std_logic;
signal un5_beamx_3_0 : std_logic;
signal un5_beamx_4 : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \beamX_RNI5457Z0Z_5\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUCZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJNZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MNZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal un5_visibley_cry_2 : std_logic;
signal un5_visibley_cry_3 : std_logic;
signal un5_visibley_cry_4 : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum\ : std_logic;
signal un5_visibley_cry_5 : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum\ : std_logic;
signal un5_visibley_cry_6 : std_logic;
signal \un5_visibley_cry_7_c_RNI1L4CZ0\ : std_logic;
signal un5_visibley_cry_7 : std_logic;
signal un5_visibley_cry_8 : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\ : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal \un4_beamylt6_cascade_\ : std_logic;
signal \un4_beamylt8_0_cascade_\ : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal \un1_beamylto9_2_cascade_\ : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal \VSync_c\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal un18_beamylt4 : std_logic;
signal \un18_beamylt4_cascade_\ : std_logic;
signal \un13_beamylt7_cascade_\ : std_logic;
signal un8_beamy_2 : std_logic;
signal un1_beamy_4 : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal un5_beamx_3 : std_logic;
signal \un8_beamylto9_1_cascade_\ : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal un5_visiblex_cry_0 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal un5_visiblex_cry_1 : std_logic;
signal un5_visiblex_cry_2 : std_logic;
signal un5_visiblex_cry_3 : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un40_sum_c5_cascade_\ : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal \un1_beamxlt10_0_cascade_\ : std_logic;
signal \HSync_c\ : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal un18_beamylto9_2 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal un1_beamx_2 : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5URZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9KZ0Z61\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02_cascade_\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8ILZ0Z1\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFRZ0Z2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6BZ0Z3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3RZ0Z3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3OZ0Z4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFEZ0Z7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7UZ0Z7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\ : std_logic;
signal \G_6_i_a4_0_0\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0_cascade_\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59\ : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0\ : std_logic;
signal un5_visibley_i : std_logic;
signal \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0\ : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal \Pixel_1_RNOZ0Z_12\ : std_logic;
signal \N_8_cascade_\ : std_logic;
signal \N_11\ : std_logic;
signal \un15_0_1_cascade_\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal un13_beamy : std_logic;
signal un4_beamy_0 : std_logic;
signal un18_beamylt10_0 : std_logic;
signal \Pixel_0_sqmuxa_0\ : std_logic;
signal \Pixel_0_sqmuxa_3\ : std_logic;
signal un1_visiblex_24 : std_logic;
signal un14lt10 : std_logic;
signal un1_visiblex_27 : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_c5_i : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un40_sum_c5 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \un5_visiblex_cry_7_c_RNIVZ0Z952\ : std_logic;
signal un5_visiblex_i_24 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \Pixel_1_RNOZ0Z_8\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PBZ0\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_i : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6\ : std_logic;
signal \bfn_12_6_0_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un54_sum_i : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2_cascade_\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\ : std_logic;
signal \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKLZ0Z62\ : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum : std_logic;
signal un1_visiblex_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PixelDebug_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    PixelDebug <= \PixelDebug_wire\;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    Pixel <= \Pixel_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    HSyncDebug <= \HSyncDebug_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__2237\,
            RESETB => \N__4336\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4866\,
            DIN => \N__4865\,
            DOUT => \N__4864\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4866\,
            PADOUT => \N__4865\,
            PADIN => \N__4864\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4082\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4857\,
            DIN => \N__4856\,
            DOUT => \N__4855\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4857\,
            PADOUT => \N__4856\,
            PADIN => \N__4855\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4848\,
            DIN => \N__4847\,
            DOUT => \N__4846\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4848\,
            PADOUT => \N__4847\,
            PADIN => \N__4846\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3481\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4839\,
            DIN => \N__4838\,
            DOUT => \N__4837\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4839\,
            PADOUT => \N__4838\,
            PADIN => \N__4837\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4069\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4830\,
            DIN => \N__4829\,
            DOUT => \N__4828\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4830\,
            PADOUT => \N__4829\,
            PADIN => \N__4828\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2831\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4821\,
            DIN => \N__4820\,
            DOUT => \N__4819\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4821\,
            PADOUT => \N__4820\,
            PADIN => \N__4819\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4812\,
            DIN => \N__4811\,
            DOUT => \N__4810\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4812\,
            PADOUT => \N__4811\,
            PADIN => \N__4810\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3482\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1051\ : InMux
    port map (
            O => \N__4793\,
            I => \N__4790\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__4790\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__4787\,
            I => \N__4784\
        );

    \I__1048\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4781\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_i
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__4778\,
            I => \N__4775\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4772\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4769\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__4760\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4751\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4751\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332\
        );

    \I__1036\ : InMux
    port map (
            O => \N__4748\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__1035\ : InMux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__4742\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__1033\ : InMux
    port map (
            O => \N__4739\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__1032\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4733\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__1030\ : InMux
    port map (
            O => \N__4730\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__1029\ : InMux
    port map (
            O => \N__4727\,
            I => \N__4723\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4720\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__4723\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__4720\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__4715\,
            I => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2_cascade_\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4706\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4706\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4706\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__4703\,
            I => \N__4699\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4694\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4694\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4694\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4686\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4681\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4681\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__4686\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__4681\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4673\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKLZ0Z62\
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__4670\,
            I => \N__4666\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4661\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4661\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__1006\ : Odrv12
    port map (
            O => \N__4658\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4652\,
            I => \N__4649\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__4649\,
            I => un1_visiblex_if_generate_plus_mult1_un61_sum_i
        );

    \I__1002\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4640\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4640\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4640\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__999\ : InMux
    port map (
            O => \N__4637\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__998\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4628\
        );

    \I__997\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4628\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4628\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PBZ0\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__994\ : InMux
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4619\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_i
        );

    \I__992\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4612\
        );

    \I__991\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4609\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__4612\,
            I => \N__4606\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4609\,
            I => \N__4603\
        );

    \I__988\ : Span4Mux_s3_h
    port map (
            O => \N__4606\,
            I => \N__4600\
        );

    \I__987\ : Span4Mux_s3_h
    port map (
            O => \N__4603\,
            I => \N__4597\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__4600\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__985\ : Odrv4
    port map (
            O => \N__4597\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum
        );

    \I__984\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4589\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03\
        );

    \I__982\ : InMux
    port map (
            O => \N__4586\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__980\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4577\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4\
        );

    \I__978\ : InMux
    port map (
            O => \N__4574\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__977\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4568\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__975\ : InMux
    port map (
            O => \N__4565\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__974\ : InMux
    port map (
            O => \N__4562\,
            I => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__4559\,
            I => \N__4555\
        );

    \I__972\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4551\
        );

    \I__971\ : InMux
    port map (
            O => \N__4555\,
            I => \N__4546\
        );

    \I__970\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4546\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4551\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4546\,
            I => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6\
        );

    \I__967\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4534\
        );

    \I__965\ : InMux
    port map (
            O => \N__4537\,
            I => \N__4531\
        );

    \I__964\ : Span4Mux_v
    port map (
            O => \N__4534\,
            I => \N__4525\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4531\,
            I => \N__4525\
        );

    \I__962\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4522\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__4525\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_c5
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4522\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_c5
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__958\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4511\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\
        );

    \I__956\ : InMux
    port map (
            O => \N__4508\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__955\ : InMux
    port map (
            O => \N__4505\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__954\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4499\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__4496\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\
        );

    \I__951\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4489\
        );

    \I__950\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4486\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4489\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4486\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__4481\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_\
        );

    \I__946\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4475\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__944\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4466\
        );

    \I__943\ : InMux
    port map (
            O => \N__4471\,
            I => \N__4466\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4466\,
            I => \N__4463\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__4463\,
            I => \un5_visiblex_cry_7_c_RNIVZ0Z952\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__4460\,
            I => \N__4457\
        );

    \I__939\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4454\,
            I => un5_visiblex_i_24
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__4451\,
            I => \N__4447\
        );

    \I__936\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4443\
        );

    \I__935\ : InMux
    port map (
            O => \N__4447\,
            I => \N__4440\
        );

    \I__934\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4437\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4432\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4432\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4437\,
            I => \N__4429\
        );

    \I__930\ : Span4Mux_s3_h
    port map (
            O => \N__4432\,
            I => \N__4426\
        );

    \I__929\ : Span4Mux_s3_h
    port map (
            O => \N__4429\,
            I => \N__4423\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__4426\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__927\ : Odrv4
    port map (
            O => \N__4423\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum
        );

    \I__926\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4412\
        );

    \I__925\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4412\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4412\,
            I => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\
        );

    \I__923\ : InMux
    port map (
            O => \N__4409\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__922\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4403\,
            I => \Pixel_1_RNOZ0Z_8\
        );

    \I__920\ : InMux
    port map (
            O => \N__4400\,
            I => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__919\ : InMux
    port map (
            O => \N__4397\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__918\ : InMux
    port map (
            O => \N__4394\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__917\ : InMux
    port map (
            O => \N__4391\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__916\ : InMux
    port map (
            O => \N__4388\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__4385\,
            I => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_\
        );

    \I__914\ : InMux
    port map (
            O => \N__4382\,
            I => \N__4376\
        );

    \I__913\ : InMux
    port map (
            O => \N__4381\,
            I => \N__4376\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__911\ : Span4Mux_s1_h
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__4370\,
            I => un1_visiblex_if_generate_plus_mult1_un54_sum
        );

    \I__909\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__4361\,
            I => un1_visiblex_if_generate_plus_mult1_un40_sum_c5_i
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__905\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4352\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0\
        );

    \I__903\ : InMux
    port map (
            O => \N__4349\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__902\ : InMux
    port map (
            O => \N__4346\,
            I => \N__4343\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4340\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__4340\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__4337\,
            I => \N__4333\
        );

    \I__898\ : IoInMux
    port map (
            O => \N__4336\,
            I => \N__4327\
        );

    \I__897\ : InMux
    port map (
            O => \N__4333\,
            I => \N__4324\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__4332\,
            I => \N__4321\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__4331\,
            I => \N__4318\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__4330\,
            I => \N__4315\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4327\,
            I => \N__4312\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4324\,
            I => \N__4309\
        );

    \I__891\ : InMux
    port map (
            O => \N__4321\,
            I => \N__4306\
        );

    \I__890\ : InMux
    port map (
            O => \N__4318\,
            I => \N__4303\
        );

    \I__889\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4300\
        );

    \I__888\ : Span4Mux_s1_v
    port map (
            O => \N__4312\,
            I => \N__4291\
        );

    \I__887\ : Span4Mux_v
    port map (
            O => \N__4309\,
            I => \N__4286\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__4306\,
            I => \N__4279\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4303\,
            I => \N__4279\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4300\,
            I => \N__4279\
        );

    \I__883\ : InMux
    port map (
            O => \N__4299\,
            I => \N__4276\
        );

    \I__882\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4271\
        );

    \I__881\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4271\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__4296\,
            I => \N__4268\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4295\,
            I => \N__4265\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__4294\,
            I => \N__4262\
        );

    \I__877\ : Span4Mux_h
    port map (
            O => \N__4291\,
            I => \N__4257\
        );

    \I__876\ : InMux
    port map (
            O => \N__4290\,
            I => \N__4252\
        );

    \I__875\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4252\
        );

    \I__874\ : Span4Mux_h
    port map (
            O => \N__4286\,
            I => \N__4243\
        );

    \I__873\ : Span4Mux_v
    port map (
            O => \N__4279\,
            I => \N__4243\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4276\,
            I => \N__4243\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4271\,
            I => \N__4243\
        );

    \I__870\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4240\
        );

    \I__869\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4235\
        );

    \I__868\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4235\
        );

    \I__867\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4232\
        );

    \I__866\ : InMux
    port map (
            O => \N__4260\,
            I => \N__4229\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__4257\,
            I => \CONSTANT_ONE_NET\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__4252\,
            I => \CONSTANT_ONE_NET\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__4243\,
            I => \CONSTANT_ONE_NET\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4240\,
            I => \CONSTANT_ONE_NET\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4235\,
            I => \CONSTANT_ONE_NET\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4232\,
            I => \CONSTANT_ONE_NET\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4229\,
            I => \CONSTANT_ONE_NET\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__4214\,
            I => \N__4211\
        );

    \I__857\ : InMux
    port map (
            O => \N__4211\,
            I => \N__4208\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4208\,
            I => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0\
        );

    \I__855\ : InMux
    port map (
            O => \N__4205\,
            I => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__854\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4198\
        );

    \I__853\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4195\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4198\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4195\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59\
        );

    \I__850\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4186\
        );

    \I__849\ : InMux
    port map (
            O => \N__4189\,
            I => \N__4183\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4186\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4183\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4178\,
            I => \N__4174\
        );

    \I__845\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4170\
        );

    \I__844\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4167\
        );

    \I__843\ : InMux
    port map (
            O => \N__4173\,
            I => \N__4164\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4170\,
            I => un5_visibley_i
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4167\,
            I => un5_visibley_i
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4164\,
            I => un5_visibley_i
        );

    \I__839\ : InMux
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4154\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__4151\,
            I => \N__4147\
        );

    \I__836\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4142\
        );

    \I__835\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4138\
        );

    \I__834\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4135\
        );

    \I__833\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4132\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4142\,
            I => \N__4129\
        );

    \I__831\ : InMux
    port map (
            O => \N__4141\,
            I => \N__4125\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4138\,
            I => \N__4118\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4135\,
            I => \N__4118\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4132\,
            I => \N__4118\
        );

    \I__827\ : Span4Mux_v
    port map (
            O => \N__4129\,
            I => \N__4115\
        );

    \I__826\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4112\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4125\,
            I => \N__4107\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__4118\,
            I => \N__4107\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__4115\,
            I => \beamYZ0Z_1\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4112\,
            I => \beamYZ0Z_1\
        );

    \I__821\ : Odrv4
    port map (
            O => \N__4107\,
            I => \beamYZ0Z_1\
        );

    \I__820\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4097\,
            I => \Pixel_1_RNOZ0Z_12\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__4094\,
            I => \N_8_cascade_\
        );

    \I__817\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4088\,
            I => \N_11\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__4085\,
            I => \un15_0_1_cascade_\
        );

    \I__814\ : IoInMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__812\ : IoSpan4Mux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__811\ : Span4Mux_s3_h
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__810\ : Span4Mux_v
    port map (
            O => \N__4070\,
            I => \N__4066\
        );

    \I__809\ : IoInMux
    port map (
            O => \N__4069\,
            I => \N__4063\
        );

    \I__808\ : Sp12to4
    port map (
            O => \N__4066\,
            I => \N__4058\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4063\,
            I => \N__4058\
        );

    \I__806\ : Odrv12
    port map (
            O => \N__4058\,
            I => \Pixel_c\
        );

    \I__805\ : ClkMux
    port map (
            O => \N__4055\,
            I => \N__4025\
        );

    \I__804\ : ClkMux
    port map (
            O => \N__4054\,
            I => \N__4025\
        );

    \I__803\ : ClkMux
    port map (
            O => \N__4053\,
            I => \N__4025\
        );

    \I__802\ : ClkMux
    port map (
            O => \N__4052\,
            I => \N__4025\
        );

    \I__801\ : ClkMux
    port map (
            O => \N__4051\,
            I => \N__4025\
        );

    \I__800\ : ClkMux
    port map (
            O => \N__4050\,
            I => \N__4025\
        );

    \I__799\ : ClkMux
    port map (
            O => \N__4049\,
            I => \N__4025\
        );

    \I__798\ : ClkMux
    port map (
            O => \N__4048\,
            I => \N__4025\
        );

    \I__797\ : ClkMux
    port map (
            O => \N__4047\,
            I => \N__4025\
        );

    \I__796\ : ClkMux
    port map (
            O => \N__4046\,
            I => \N__4025\
        );

    \I__795\ : GlobalMux
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__794\ : gio2CtrlBuf
    port map (
            O => \N__4022\,
            I => \PixelClock_g\
        );

    \I__793\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4016\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4016\,
            I => un13_beamy
        );

    \I__791\ : InMux
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4010\,
            I => un4_beamy_0
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__4007\,
            I => \N__4004\
        );

    \I__788\ : InMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__3998\,
            I => un18_beamylt10_0
        );

    \I__785\ : InMux
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__783\ : Odrv4
    port map (
            O => \N__3989\,
            I => \Pixel_0_sqmuxa_0\
        );

    \I__782\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3983\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3983\,
            I => \Pixel_0_sqmuxa_3\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__779\ : InMux
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__3974\,
            I => \N__3971\
        );

    \I__777\ : Span4Mux_s3_h
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__3968\,
            I => un1_visiblex_24
        );

    \I__775\ : InMux
    port map (
            O => \N__3965\,
            I => \N__3962\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__3962\,
            I => \N__3959\
        );

    \I__773\ : Odrv12
    port map (
            O => \N__3959\,
            I => un14lt10
        );

    \I__772\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3953\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3953\,
            I => \N__3950\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__3950\,
            I => un1_visiblex_27
        );

    \I__769\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3943\
        );

    \I__768\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3940\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__3943\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3940\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__3935\,
            I => \N__3932\
        );

    \I__764\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3929\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\
        );

    \I__762\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3923\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__3923\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\
        );

    \I__760\ : InMux
    port map (
            O => \N__3920\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__3917\,
            I => \N__3914\
        );

    \I__758\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3911\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3OZ0Z4\
        );

    \I__756\ : InMux
    port map (
            O => \N__3908\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\
        );

    \I__755\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3902\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFEZ0Z7\
        );

    \I__753\ : InMux
    port map (
            O => \N__3899\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\
        );

    \I__752\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3893\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7UZ0Z7\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__3890\,
            I => \N__3885\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__3889\,
            I => \N__3881\
        );

    \I__748\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3877\
        );

    \I__747\ : InMux
    port map (
            O => \N__3885\,
            I => \N__3868\
        );

    \I__746\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3868\
        );

    \I__745\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3868\
        );

    \I__744\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3868\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__3877\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3868\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__740\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3857\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\
        );

    \I__738\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__3851\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\
        );

    \I__736\ : InMux
    port map (
            O => \N__3848\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\
        );

    \I__735\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3842\,
            I => \G_6_i_a4_0_0\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__3839\,
            I => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0_cascade_\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__3836\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4_cascade_\
        );

    \I__731\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3829\
        );

    \I__730\ : InMux
    port map (
            O => \N__3832\,
            I => \N__3826\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3829\,
            I => \N__3823\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3826\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__727\ : Odrv4
    port map (
            O => \N__3823\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__3818\,
            I => \N__3815\
        );

    \I__725\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3812\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3812\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\
        );

    \I__723\ : InMux
    port map (
            O => \N__3809\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\
        );

    \I__722\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3803\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3803\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFRZ0Z2\
        );

    \I__720\ : InMux
    port map (
            O => \N__3800\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__3797\,
            I => \N__3793\
        );

    \I__718\ : InMux
    port map (
            O => \N__3796\,
            I => \N__3784\
        );

    \I__717\ : InMux
    port map (
            O => \N__3793\,
            I => \N__3784\
        );

    \I__716\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3784\
        );

    \I__715\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3781\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3784\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__3781\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__3776\,
            I => \N__3773\
        );

    \I__711\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3770\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6BZ0Z3\
        );

    \I__709\ : InMux
    port map (
            O => \N__3767\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\
        );

    \I__708\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3761\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__3761\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3RZ0Z3\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__3758\,
            I => \N__3755\
        );

    \I__705\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3752\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__3752\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\
        );

    \I__703\ : InMux
    port map (
            O => \N__3749\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\
        );

    \I__702\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3743\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\
        );

    \I__700\ : InMux
    port map (
            O => \N__3740\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__3737\,
            I => \N__3733\
        );

    \I__698\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3728\
        );

    \I__697\ : InMux
    port map (
            O => \N__3733\,
            I => \N__3728\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3728\,
            I => \un1_beamY_if_generate_plus_mult1_un68_sum\
        );

    \I__695\ : InMux
    port map (
            O => \N__3725\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\
        );

    \I__694\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3719\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\
        );

    \I__692\ : InMux
    port map (
            O => \N__3716\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__3713\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02_cascade_\
        );

    \I__690\ : InMux
    port map (
            O => \N__3710\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\
        );

    \I__689\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3704\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\
        );

    \I__687\ : InMux
    port map (
            O => \N__3701\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__3698\,
            I => \N__3694\
        );

    \I__685\ : InMux
    port map (
            O => \N__3697\,
            I => \N__3685\
        );

    \I__684\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3685\
        );

    \I__683\ : InMux
    port map (
            O => \N__3693\,
            I => \N__3685\
        );

    \I__682\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3682\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3685\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3682\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__678\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3671\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\
        );

    \I__676\ : InMux
    port map (
            O => \N__3668\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\
        );

    \I__675\ : InMux
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3662\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8ILZ0Z1\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__672\ : InMux
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3653\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\
        );

    \I__670\ : InMux
    port map (
            O => \N__3650\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\
        );

    \I__669\ : InMux
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__3644\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\
        );

    \I__667\ : InMux
    port map (
            O => \N__3641\,
            I => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__3638\,
            I => \N__3635\
        );

    \I__665\ : InMux
    port map (
            O => \N__3635\,
            I => \N__3628\
        );

    \I__664\ : InMux
    port map (
            O => \N__3634\,
            I => \N__3623\
        );

    \I__663\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3623\
        );

    \I__662\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3619\
        );

    \I__661\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3616\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3628\,
            I => \N__3613\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3623\,
            I => \N__3610\
        );

    \I__658\ : InMux
    port map (
            O => \N__3622\,
            I => \N__3607\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__3619\,
            I => \beamXZ0Z_5\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3616\,
            I => \beamXZ0Z_5\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__3613\,
            I => \beamXZ0Z_5\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__3610\,
            I => \beamXZ0Z_5\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3607\,
            I => \beamXZ0Z_5\
        );

    \I__652\ : InMux
    port map (
            O => \N__3596\,
            I => \N__3589\
        );

    \I__651\ : InMux
    port map (
            O => \N__3595\,
            I => \N__3584\
        );

    \I__650\ : InMux
    port map (
            O => \N__3594\,
            I => \N__3584\
        );

    \I__649\ : InMux
    port map (
            O => \N__3593\,
            I => \N__3580\
        );

    \I__648\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3577\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3589\,
            I => \N__3574\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3584\,
            I => \N__3571\
        );

    \I__645\ : InMux
    port map (
            O => \N__3583\,
            I => \N__3568\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3580\,
            I => \beamXZ0Z_4\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3577\,
            I => \beamXZ0Z_4\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__3574\,
            I => \beamXZ0Z_4\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__3571\,
            I => \beamXZ0Z_4\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3568\,
            I => \beamXZ0Z_4\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3557\,
            I => \N__3553\
        );

    \I__638\ : InMux
    port map (
            O => \N__3556\,
            I => \N__3548\
        );

    \I__637\ : InMux
    port map (
            O => \N__3553\,
            I => \N__3545\
        );

    \I__636\ : InMux
    port map (
            O => \N__3552\,
            I => \N__3541\
        );

    \I__635\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3538\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3548\,
            I => \N__3533\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3545\,
            I => \N__3533\
        );

    \I__632\ : InMux
    port map (
            O => \N__3544\,
            I => \N__3530\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3541\,
            I => \beamXZ0Z_3\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3538\,
            I => \beamXZ0Z_3\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__3533\,
            I => \beamXZ0Z_3\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3530\,
            I => \beamXZ0Z_3\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__3521\,
            I => \N__3516\
        );

    \I__626\ : InMux
    port map (
            O => \N__3520\,
            I => \N__3511\
        );

    \I__625\ : InMux
    port map (
            O => \N__3519\,
            I => \N__3511\
        );

    \I__624\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3508\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3511\,
            I => \N__3501\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__3508\,
            I => \N__3501\
        );

    \I__621\ : InMux
    port map (
            O => \N__3507\,
            I => \N__3498\
        );

    \I__620\ : InMux
    port map (
            O => \N__3506\,
            I => \N__3495\
        );

    \I__619\ : Span4Mux_h
    port map (
            O => \N__3501\,
            I => \N__3492\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3498\,
            I => \beamXZ0Z_10\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__3495\,
            I => \beamXZ0Z_10\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__3492\,
            I => \beamXZ0Z_10\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__3485\,
            I => \un1_beamxlt10_0_cascade_\
        );

    \I__614\ : IoInMux
    port map (
            O => \N__3482\,
            I => \N__3478\
        );

    \I__613\ : IoInMux
    port map (
            O => \N__3481\,
            I => \N__3475\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3478\,
            I => \N__3472\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3475\,
            I => \N__3469\
        );

    \I__610\ : Span12Mux_s9_v
    port map (
            O => \N__3472\,
            I => \N__3466\
        );

    \I__609\ : Span4Mux_s2_v
    port map (
            O => \N__3469\,
            I => \N__3463\
        );

    \I__608\ : Odrv12
    port map (
            O => \N__3466\,
            I => \HSync_c\
        );

    \I__607\ : Odrv4
    port map (
            O => \N__3463\,
            I => \HSync_c\
        );

    \I__606\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3454\
        );

    \I__605\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3450\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3454\,
            I => \N__3444\
        );

    \I__603\ : InMux
    port map (
            O => \N__3453\,
            I => \N__3441\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3450\,
            I => \N__3438\
        );

    \I__601\ : InMux
    port map (
            O => \N__3449\,
            I => \N__3433\
        );

    \I__600\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3433\
        );

    \I__599\ : InMux
    port map (
            O => \N__3447\,
            I => \N__3430\
        );

    \I__598\ : Odrv4
    port map (
            O => \N__3444\,
            I => \beamXZ0Z_7\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3441\,
            I => \beamXZ0Z_7\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__3438\,
            I => \beamXZ0Z_7\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3433\,
            I => \beamXZ0Z_7\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3430\,
            I => \beamXZ0Z_7\
        );

    \I__593\ : InMux
    port map (
            O => \N__3419\,
            I => \N__3415\
        );

    \I__592\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3412\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3415\,
            I => \N__3405\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3412\,
            I => \N__3405\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__3411\,
            I => \N__3402\
        );

    \I__588\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3397\
        );

    \I__587\ : Span4Mux_h
    port map (
            O => \N__3405\,
            I => \N__3394\
        );

    \I__586\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3389\
        );

    \I__585\ : InMux
    port map (
            O => \N__3401\,
            I => \N__3389\
        );

    \I__584\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3386\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3397\,
            I => \beamXZ0Z_6\
        );

    \I__582\ : Odrv4
    port map (
            O => \N__3394\,
            I => \beamXZ0Z_6\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3389\,
            I => \beamXZ0Z_6\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3386\,
            I => \beamXZ0Z_6\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__578\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3371\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__3368\,
            I => un18_beamylto9_2
        );

    \I__575\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3359\
        );

    \I__574\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3356\
        );

    \I__573\ : InMux
    port map (
            O => \N__3363\,
            I => \N__3351\
        );

    \I__572\ : InMux
    port map (
            O => \N__3362\,
            I => \N__3351\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3359\,
            I => \beamXZ0Z_8\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3356\,
            I => \beamXZ0Z_8\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3351\,
            I => \beamXZ0Z_8\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__3344\,
            I => \N__3340\
        );

    \I__567\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3335\
        );

    \I__566\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3328\
        );

    \I__565\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3328\
        );

    \I__564\ : InMux
    port map (
            O => \N__3338\,
            I => \N__3328\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3335\,
            I => \beamXZ0Z_9\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3328\,
            I => \beamXZ0Z_9\
        );

    \I__561\ : InMux
    port map (
            O => \N__3323\,
            I => \N__3318\
        );

    \I__560\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3315\
        );

    \I__559\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3312\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3318\,
            I => \N__3307\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3315\,
            I => \N__3307\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3312\,
            I => un1_beamx_2
        );

    \I__555\ : Odrv4
    port map (
            O => \N__3307\,
            I => un1_beamx_2
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__553\ : InMux
    port map (
            O => \N__3299\,
            I => \N__3296\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3296\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\
        );

    \I__551\ : InMux
    port map (
            O => \N__3293\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\
        );

    \I__550\ : InMux
    port map (
            O => \N__3290\,
            I => \N__3287\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3287\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\
        );

    \I__548\ : InMux
    port map (
            O => \N__3284\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__3281\,
            I => \N__3277\
        );

    \I__546\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3268\
        );

    \I__545\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3268\
        );

    \I__544\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3268\
        );

    \I__543\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3265\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3268\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3265\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__3260\,
            I => \N__3257\
        );

    \I__539\ : InMux
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3254\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5URZ0\
        );

    \I__537\ : InMux
    port map (
            O => \N__3251\,
            I => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\
        );

    \I__536\ : InMux
    port map (
            O => \N__3248\,
            I => \N__3245\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__3245\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9KZ0Z61\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__3242\,
            I => \N__3239\
        );

    \I__533\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3236\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\
        );

    \I__531\ : InMux
    port map (
            O => \N__3233\,
            I => \N__3227\
        );

    \I__530\ : InMux
    port map (
            O => \N__3232\,
            I => \N__3224\
        );

    \I__529\ : InMux
    port map (
            O => \N__3231\,
            I => \N__3221\
        );

    \I__528\ : InMux
    port map (
            O => \N__3230\,
            I => \N__3218\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3227\,
            I => \N__3213\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3224\,
            I => \N__3213\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3221\,
            I => \N__3210\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3218\,
            I => \beamXZ0Z_2\
        );

    \I__523\ : Odrv4
    port map (
            O => \N__3213\,
            I => \beamXZ0Z_2\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__3210\,
            I => \beamXZ0Z_2\
        );

    \I__521\ : InMux
    port map (
            O => \N__3203\,
            I => un5_visiblex_cry_2
        );

    \I__520\ : InMux
    port map (
            O => \N__3200\,
            I => un5_visiblex_cry_3
        );

    \I__519\ : InMux
    port map (
            O => \N__3197\,
            I => un5_visiblex_cry_4
        );

    \I__518\ : InMux
    port map (
            O => \N__3194\,
            I => un5_visiblex_cry_5
        );

    \I__517\ : InMux
    port map (
            O => \N__3191\,
            I => un5_visiblex_cry_6
        );

    \I__516\ : InMux
    port map (
            O => \N__3188\,
            I => \bfn_8_7_0_\
        );

    \I__515\ : InMux
    port map (
            O => \N__3185\,
            I => un5_visiblex_cry_8
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__3182\,
            I => \un1_visiblex_if_generate_plus_mult1_un40_sum_c5_cascade_\
        );

    \I__513\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3176\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3176\,
            I => un18_beamylt4
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3173\,
            I => \un18_beamylt4_cascade_\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__3170\,
            I => \un13_beamylt7_cascade_\
        );

    \I__509\ : InMux
    port map (
            O => \N__3167\,
            I => \N__3164\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3164\,
            I => \N__3160\
        );

    \I__507\ : InMux
    port map (
            O => \N__3163\,
            I => \N__3157\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__3160\,
            I => un8_beamy_2
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3157\,
            I => un8_beamy_2
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3152\,
            I => \N__3147\
        );

    \I__503\ : InMux
    port map (
            O => \N__3151\,
            I => \N__3144\
        );

    \I__502\ : InMux
    port map (
            O => \N__3150\,
            I => \N__3141\
        );

    \I__501\ : InMux
    port map (
            O => \N__3147\,
            I => \N__3138\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3144\,
            I => \N__3135\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3141\,
            I => un1_beamy_4
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3138\,
            I => un1_beamy_4
        );

    \I__497\ : Odrv4
    port map (
            O => \N__3135\,
            I => un1_beamy_4
        );

    \I__496\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3124\
        );

    \I__495\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3121\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3124\,
            I => \N__3112\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3121\,
            I => \N__3112\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__3120\,
            I => \N__3109\
        );

    \I__491\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3106\
        );

    \I__490\ : InMux
    port map (
            O => \N__3118\,
            I => \N__3103\
        );

    \I__489\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3100\
        );

    \I__488\ : Span4Mux_v
    port map (
            O => \N__3112\,
            I => \N__3097\
        );

    \I__487\ : InMux
    port map (
            O => \N__3109\,
            I => \N__3094\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3106\,
            I => \beamYZ0Z_7\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3103\,
            I => \beamYZ0Z_7\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3100\,
            I => \beamYZ0Z_7\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3097\,
            I => \beamYZ0Z_7\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3094\,
            I => \beamYZ0Z_7\
        );

    \I__481\ : InMux
    port map (
            O => \N__3083\,
            I => \N__3073\
        );

    \I__480\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3073\
        );

    \I__479\ : InMux
    port map (
            O => \N__3081\,
            I => \N__3063\
        );

    \I__478\ : InMux
    port map (
            O => \N__3080\,
            I => \N__3063\
        );

    \I__477\ : InMux
    port map (
            O => \N__3079\,
            I => \N__3063\
        );

    \I__476\ : InMux
    port map (
            O => \N__3078\,
            I => \N__3063\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__3073\,
            I => \N__3060\
        );

    \I__474\ : InMux
    port map (
            O => \N__3072\,
            I => \N__3057\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3063\,
            I => un5_beamx_3
        );

    \I__472\ : Odrv4
    port map (
            O => \N__3060\,
            I => un5_beamx_3
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3057\,
            I => un5_beamx_3
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__3050\,
            I => \un8_beamylto9_1_cascade_\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__3047\,
            I => \N__3043\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3046\,
            I => \N__3035\
        );

    \I__467\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3032\
        );

    \I__466\ : InMux
    port map (
            O => \N__3042\,
            I => \N__3029\
        );

    \I__465\ : InMux
    port map (
            O => \N__3041\,
            I => \N__3026\
        );

    \I__464\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3019\
        );

    \I__463\ : InMux
    port map (
            O => \N__3039\,
            I => \N__3019\
        );

    \I__462\ : InMux
    port map (
            O => \N__3038\,
            I => \N__3019\
        );

    \I__461\ : InMux
    port map (
            O => \N__3035\,
            I => \N__3016\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3032\,
            I => \beamYZ0Z_2\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3029\,
            I => \beamYZ0Z_2\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3026\,
            I => \beamYZ0Z_2\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3019\,
            I => \beamYZ0Z_2\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3016\,
            I => \beamYZ0Z_2\
        );

    \I__455\ : InMux
    port map (
            O => \N__3005\,
            I => \N__3002\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__3002\,
            I => \N__2994\
        );

    \I__453\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2989\
        );

    \I__452\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2989\
        );

    \I__451\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2986\
        );

    \I__450\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2981\
        );

    \I__449\ : InMux
    port map (
            O => \N__2997\,
            I => \N__2981\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__2994\,
            I => \beamXZ0Z_0\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__2989\,
            I => \beamXZ0Z_0\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2986\,
            I => \beamXZ0Z_0\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2981\,
            I => \beamXZ0Z_0\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__2972\,
            I => \N__2969\
        );

    \I__443\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2963\
        );

    \I__442\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2960\
        );

    \I__441\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2957\
        );

    \I__440\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2954\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2963\,
            I => \beamXZ0Z_1\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2960\,
            I => \beamXZ0Z_1\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2957\,
            I => \beamXZ0Z_1\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2954\,
            I => \beamXZ0Z_1\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__2945\,
            I => \N__2939\
        );

    \I__434\ : InMux
    port map (
            O => \N__2944\,
            I => \N__2936\
        );

    \I__433\ : InMux
    port map (
            O => \N__2943\,
            I => \N__2933\
        );

    \I__432\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2930\
        );

    \I__431\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2927\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2936\,
            I => \beamYZ0Z_6\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2933\,
            I => \beamYZ0Z_6\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2930\,
            I => \beamYZ0Z_6\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__2927\,
            I => \beamYZ0Z_6\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__2918\,
            I => \N__2912\
        );

    \I__425\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2909\
        );

    \I__424\ : InMux
    port map (
            O => \N__2916\,
            I => \N__2904\
        );

    \I__423\ : InMux
    port map (
            O => \N__2915\,
            I => \N__2904\
        );

    \I__422\ : InMux
    port map (
            O => \N__2912\,
            I => \N__2901\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2909\,
            I => \beamYZ0Z_5\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__2904\,
            I => \beamYZ0Z_5\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2901\,
            I => \beamYZ0Z_5\
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__2894\,
            I => \un4_beamylt6_cascade_\
        );

    \I__417\ : CascadeMux
    port map (
            O => \N__2891\,
            I => \un4_beamylt8_0_cascade_\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__2888\,
            I => \N__2881\
        );

    \I__415\ : InMux
    port map (
            O => \N__2887\,
            I => \N__2878\
        );

    \I__414\ : InMux
    port map (
            O => \N__2886\,
            I => \N__2871\
        );

    \I__413\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2871\
        );

    \I__412\ : InMux
    port map (
            O => \N__2884\,
            I => \N__2871\
        );

    \I__411\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2868\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__2878\,
            I => \beamYZ0Z_3\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2871\,
            I => \beamYZ0Z_3\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2868\,
            I => \beamYZ0Z_3\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__2861\,
            I => \un1_beamylto9_2_cascade_\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__2858\,
            I => \N__2851\
        );

    \I__405\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2848\
        );

    \I__404\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2841\
        );

    \I__403\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2841\
        );

    \I__402\ : InMux
    port map (
            O => \N__2854\,
            I => \N__2841\
        );

    \I__401\ : InMux
    port map (
            O => \N__2851\,
            I => \N__2838\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2848\,
            I => \beamYZ0Z_4\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2841\,
            I => \beamYZ0Z_4\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__2838\,
            I => \beamYZ0Z_4\
        );

    \I__397\ : IoInMux
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2828\,
            I => \N__2825\
        );

    \I__395\ : IoSpan4Mux
    port map (
            O => \N__2825\,
            I => \N__2822\
        );

    \I__394\ : Sp12to4
    port map (
            O => \N__2822\,
            I => \N__2818\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__2821\,
            I => \N__2815\
        );

    \I__392\ : Span12Mux_v
    port map (
            O => \N__2818\,
            I => \N__2812\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2815\,
            I => \N__2809\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__2812\,
            I => \VSync_c\
        );

    \I__389\ : Odrv12
    port map (
            O => \N__2809\,
            I => \VSync_c\
        );

    \I__388\ : InMux
    port map (
            O => \N__2804\,
            I => \N__2796\
        );

    \I__387\ : InMux
    port map (
            O => \N__2803\,
            I => \N__2796\
        );

    \I__386\ : InMux
    port map (
            O => \N__2802\,
            I => \N__2793\
        );

    \I__385\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2789\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__2796\,
            I => \N__2784\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2793\,
            I => \N__2784\
        );

    \I__382\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2781\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__2789\,
            I => \beamYZ0Z_9\
        );

    \I__380\ : Odrv4
    port map (
            O => \N__2784\,
            I => \beamYZ0Z_9\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2781\,
            I => \beamYZ0Z_9\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__2774\,
            I => \N__2767\
        );

    \I__377\ : InMux
    port map (
            O => \N__2773\,
            I => \N__2764\
        );

    \I__376\ : InMux
    port map (
            O => \N__2772\,
            I => \N__2761\
        );

    \I__375\ : InMux
    port map (
            O => \N__2771\,
            I => \N__2758\
        );

    \I__374\ : InMux
    port map (
            O => \N__2770\,
            I => \N__2755\
        );

    \I__373\ : InMux
    port map (
            O => \N__2767\,
            I => \N__2752\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__2764\,
            I => \beamYZ0Z_8\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2761\,
            I => \beamYZ0Z_8\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2758\,
            I => \beamYZ0Z_8\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2755\,
            I => \beamYZ0Z_8\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2752\,
            I => \beamYZ0Z_8\
        );

    \I__367\ : InMux
    port map (
            O => \N__2741\,
            I => un5_visibley_cry_2
        );

    \I__366\ : InMux
    port map (
            O => \N__2738\,
            I => un5_visibley_cry_3
        );

    \I__365\ : InMux
    port map (
            O => \N__2735\,
            I => un5_visibley_cry_4
        );

    \I__364\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2728\
        );

    \I__363\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2725\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2728\,
            I => \N__2722\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2725\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__2722\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum\
        );

    \I__359\ : InMux
    port map (
            O => \N__2717\,
            I => un5_visibley_cry_5
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__357\ : InMux
    port map (
            O => \N__2711\,
            I => \N__2707\
        );

    \I__356\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2704\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2707\,
            I => \N__2701\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__2704\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__353\ : Odrv4
    port map (
            O => \N__2701\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum\
        );

    \I__352\ : InMux
    port map (
            O => \N__2696\,
            I => un5_visibley_cry_6
        );

    \I__351\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2687\
        );

    \I__350\ : InMux
    port map (
            O => \N__2692\,
            I => \N__2687\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2687\,
            I => \un5_visibley_cry_7_c_RNI1L4CZ0\
        );

    \I__348\ : InMux
    port map (
            O => \N__2684\,
            I => un5_visibley_cry_7
        );

    \I__347\ : InMux
    port map (
            O => \N__2681\,
            I => un5_visibley_cry_8
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__2678\,
            I => \N__2675\
        );

    \I__345\ : InMux
    port map (
            O => \N__2675\,
            I => \N__2669\
        );

    \I__344\ : InMux
    port map (
            O => \N__2674\,
            I => \N__2669\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2669\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\
        );

    \I__342\ : CEMux
    port map (
            O => \N__2666\,
            I => \N__2661\
        );

    \I__341\ : InMux
    port map (
            O => \N__2665\,
            I => \N__2656\
        );

    \I__340\ : InMux
    port map (
            O => \N__2664\,
            I => \N__2653\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2661\,
            I => \N__2650\
        );

    \I__338\ : CEMux
    port map (
            O => \N__2660\,
            I => \N__2647\
        );

    \I__337\ : CEMux
    port map (
            O => \N__2659\,
            I => \N__2643\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__2656\,
            I => \N__2634\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2653\,
            I => \N__2634\
        );

    \I__334\ : Span4Mux_v
    port map (
            O => \N__2650\,
            I => \N__2634\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2647\,
            I => \N__2634\
        );

    \I__332\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2631\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2643\,
            I => \N__2626\
        );

    \I__330\ : Span4Mux_v
    port map (
            O => \N__2634\,
            I => \N__2626\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2631\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__328\ : Odrv4
    port map (
            O => \N__2626\,
            I => \beamX_RNI5457Z0Z_5\
        );

    \I__327\ : InMux
    port map (
            O => \N__2621\,
            I => un8_beamx_cry_9
        );

    \I__326\ : InMux
    port map (
            O => \N__2618\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\
        );

    \I__325\ : CascadeMux
    port map (
            O => \N__2615\,
            I => \N__2612\
        );

    \I__324\ : InMux
    port map (
            O => \N__2612\,
            I => \N__2609\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2609\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUCZ0\
        );

    \I__322\ : InMux
    port map (
            O => \N__2606\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\
        );

    \I__321\ : InMux
    port map (
            O => \N__2603\,
            I => \N__2600\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2600\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJNZ0\
        );

    \I__319\ : InMux
    port map (
            O => \N__2597\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\
        );

    \I__318\ : InMux
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__2591\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MNZ0\
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__2588\,
            I => \N__2585\
        );

    \I__315\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2582\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\
        );

    \I__313\ : InMux
    port map (
            O => \N__2579\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\
        );

    \I__312\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2573\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__310\ : CascadeMux
    port map (
            O => \N__2570\,
            I => \N__2565\
        );

    \I__309\ : InMux
    port map (
            O => \N__2569\,
            I => \N__2562\
        );

    \I__308\ : InMux
    port map (
            O => \N__2568\,
            I => \N__2559\
        );

    \I__307\ : InMux
    port map (
            O => \N__2565\,
            I => \N__2556\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2562\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__2559\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2556\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\
        );

    \I__303\ : CascadeMux
    port map (
            O => \N__2549\,
            I => \N__2544\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__2548\,
            I => \N__2541\
        );

    \I__301\ : CascadeMux
    port map (
            O => \N__2547\,
            I => \N__2537\
        );

    \I__300\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2528\
        );

    \I__299\ : InMux
    port map (
            O => \N__2541\,
            I => \N__2528\
        );

    \I__298\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2528\
        );

    \I__297\ : InMux
    port map (
            O => \N__2537\,
            I => \N__2528\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2528\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\
        );

    \I__295\ : InMux
    port map (
            O => \N__2525\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\
        );

    \I__294\ : CascadeMux
    port map (
            O => \N__2522\,
            I => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\
        );

    \I__293\ : InMux
    port map (
            O => \N__2519\,
            I => \N__2516\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2516\,
            I => \N__2513\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__2513\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\
        );

    \I__290\ : InMux
    port map (
            O => \N__2510\,
            I => un8_beamx_cry_1
        );

    \I__289\ : InMux
    port map (
            O => \N__2507\,
            I => un8_beamx_cry_2
        );

    \I__288\ : InMux
    port map (
            O => \N__2504\,
            I => un8_beamx_cry_3
        );

    \I__287\ : InMux
    port map (
            O => \N__2501\,
            I => un8_beamx_cry_4
        );

    \I__286\ : InMux
    port map (
            O => \N__2498\,
            I => un8_beamx_cry_5
        );

    \I__285\ : InMux
    port map (
            O => \N__2495\,
            I => un8_beamx_cry_6
        );

    \I__284\ : InMux
    port map (
            O => \N__2492\,
            I => un8_beamx_cry_7
        );

    \I__283\ : InMux
    port map (
            O => \N__2489\,
            I => \bfn_7_8_0_\
        );

    \I__282\ : InMux
    port map (
            O => \N__2486\,
            I => \bfn_7_5_0_\
        );

    \I__281\ : InMux
    port map (
            O => \N__2483\,
            I => \N__2480\
        );

    \I__280\ : LocalMux
    port map (
            O => \N__2480\,
            I => \N__2477\
        );

    \I__279\ : Odrv4
    port map (
            O => \N__2477\,
            I => \beamY_RNO_0Z0Z_9\
        );

    \I__278\ : CascadeMux
    port map (
            O => \N__2474\,
            I => \un3_beamx_5_cascade_\
        );

    \I__277\ : InMux
    port map (
            O => \N__2471\,
            I => \N__2468\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2468\,
            I => un3_beamx_7
        );

    \I__275\ : InMux
    port map (
            O => \N__2465\,
            I => \N__2462\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2462\,
            I => \beamY_RNO_0Z0Z_1\
        );

    \I__273\ : CascadeMux
    port map (
            O => \N__2459\,
            I => \N__2456\
        );

    \I__272\ : InMux
    port map (
            O => \N__2456\,
            I => \N__2444\
        );

    \I__271\ : InMux
    port map (
            O => \N__2455\,
            I => \N__2444\
        );

    \I__270\ : InMux
    port map (
            O => \N__2454\,
            I => \N__2444\
        );

    \I__269\ : InMux
    port map (
            O => \N__2453\,
            I => \N__2444\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2444\,
            I => \N__2439\
        );

    \I__267\ : InMux
    port map (
            O => \N__2443\,
            I => \N__2434\
        );

    \I__266\ : InMux
    port map (
            O => \N__2442\,
            I => \N__2434\
        );

    \I__265\ : Odrv4
    port map (
            O => \N__2439\,
            I => un5_beamx_3_0
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2434\,
            I => un5_beamx_3_0
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__2429\,
            I => \N__2423\
        );

    \I__262\ : InMux
    port map (
            O => \N__2428\,
            I => \N__2413\
        );

    \I__261\ : InMux
    port map (
            O => \N__2427\,
            I => \N__2413\
        );

    \I__260\ : InMux
    port map (
            O => \N__2426\,
            I => \N__2413\
        );

    \I__259\ : InMux
    port map (
            O => \N__2423\,
            I => \N__2413\
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__2422\,
            I => \N__2410\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2413\,
            I => \N__2406\
        );

    \I__256\ : InMux
    port map (
            O => \N__2410\,
            I => \N__2401\
        );

    \I__255\ : InMux
    port map (
            O => \N__2409\,
            I => \N__2401\
        );

    \I__254\ : Odrv4
    port map (
            O => \N__2406\,
            I => un5_beamx_4
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2401\,
            I => un5_beamx_4
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__2396\,
            I => \N__2392\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__2395\,
            I => \N__2389\
        );

    \I__250\ : InMux
    port map (
            O => \N__2392\,
            I => \N__2384\
        );

    \I__249\ : InMux
    port map (
            O => \N__2389\,
            I => \N__2381\
        );

    \I__248\ : InMux
    port map (
            O => \N__2388\,
            I => \N__2378\
        );

    \I__247\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2375\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2384\,
            I => \N__2372\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2381\,
            I => \beamYZ0Z_0\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__2378\,
            I => \beamYZ0Z_0\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2375\,
            I => \beamYZ0Z_0\
        );

    \I__242\ : Odrv4
    port map (
            O => \N__2372\,
            I => \beamYZ0Z_0\
        );

    \I__241\ : InMux
    port map (
            O => \N__2363\,
            I => un21_beamy_cry_1
        );

    \I__240\ : InMux
    port map (
            O => \N__2360\,
            I => \N__2357\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2357\,
            I => \beamY_RNO_0Z0Z_3\
        );

    \I__238\ : InMux
    port map (
            O => \N__2354\,
            I => un21_beamy_cry_2
        );

    \I__237\ : CascadeMux
    port map (
            O => \N__2351\,
            I => \N__2348\
        );

    \I__236\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2345\,
            I => \beamY_RNO_0Z0Z_4\
        );

    \I__234\ : InMux
    port map (
            O => \N__2342\,
            I => un21_beamy_cry_3
        );

    \I__233\ : InMux
    port map (
            O => \N__2339\,
            I => un21_beamy_cry_4
        );

    \I__232\ : InMux
    port map (
            O => \N__2336\,
            I => un21_beamy_cry_5
        );

    \I__231\ : CascadeMux
    port map (
            O => \N__2333\,
            I => \N__2330\
        );

    \I__230\ : InMux
    port map (
            O => \N__2330\,
            I => \N__2327\
        );

    \I__229\ : LocalMux
    port map (
            O => \N__2327\,
            I => \beamY_RNO_0Z0Z_7\
        );

    \I__228\ : InMux
    port map (
            O => \N__2324\,
            I => un21_beamy_cry_6
        );

    \I__227\ : InMux
    port map (
            O => \N__2321\,
            I => un21_beamy_cry_7
        );

    \I__226\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2315\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2315\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPMZ0\
        );

    \I__224\ : InMux
    port map (
            O => \N__2312\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\
        );

    \I__223\ : InMux
    port map (
            O => \N__2309\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\
        );

    \I__222\ : InMux
    port map (
            O => \N__2306\,
            I => \N__2303\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2303\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__2300\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\
        );

    \I__219\ : CascadeMux
    port map (
            O => \N__2297\,
            I => \N__2294\
        );

    \I__218\ : InMux
    port map (
            O => \N__2294\,
            I => \N__2291\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2291\,
            I => \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\
        );

    \I__216\ : InMux
    port map (
            O => \N__2288\,
            I => \N__2285\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__2285\,
            I => \un5_visibley_cry_7_c_RNI1L4CZ0Z_0\
        );

    \I__214\ : InMux
    port map (
            O => \N__2282\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\
        );

    \I__213\ : InMux
    port map (
            O => \N__2279\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\
        );

    \I__212\ : InMux
    port map (
            O => \N__2276\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\
        );

    \I__211\ : InMux
    port map (
            O => \N__2273\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\
        );

    \I__210\ : InMux
    port map (
            O => \N__2270\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\
        );

    \I__209\ : CascadeMux
    port map (
            O => \N__2267\,
            I => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\
        );

    \I__208\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2261\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2261\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOMZ0\
        );

    \I__206\ : InMux
    port map (
            O => \N__2258\,
            I => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\
        );

    \I__205\ : IoInMux
    port map (
            O => \N__2255\,
            I => \N__2252\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2252\,
            I => \N__2249\
        );

    \I__203\ : Span4Mux_s1_h
    port map (
            O => \N__2249\,
            I => \N__2246\
        );

    \I__202\ : Span4Mux_h
    port map (
            O => \N__2246\,
            I => \N__2243\
        );

    \I__201\ : Sp12to4
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__200\ : Odrv12
    port map (
            O => \N__2240\,
            I => \Clock50MHz.PixelClock\
        );

    \I__199\ : IoInMux
    port map (
            O => \N__2237\,
            I => \N__2234\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__2234\,
            I => \N__2231\
        );

    \I__197\ : IoSpan4Mux
    port map (
            O => \N__2231\,
            I => \N__2228\
        );

    \I__196\ : Odrv4
    port map (
            O => \N__2228\,
            I => \Clock12MHz_c\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_cry_7,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un21_beamy_cry_8,
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_12_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_6_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_7_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_1_0_\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2255\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \beamY_RNO_0_1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2388\,
            in2 => \_gnd_net_\,
            in3 => \N__4128\,
            lcout => \beamY_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2714\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_1_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUC_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2288\,
            in2 => \N__4294\,
            in3 => \N__2282\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNIOQUCZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJN_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2264\,
            in2 => \N__4296\,
            in3 => \N__2279\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSJNZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MN_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2318\,
            in2 => \N__4295\,
            in3 => \N__2276\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIM0MNZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2570\,
            in3 => \N__2273\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2306\,
            in2 => \_gnd_net_\,
            in3 => \N__2270\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_0_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2267\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2692\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOM_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4260\,
            in2 => \N__2297\,
            in3 => \N__2258\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNISKOMZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPM_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4261\,
            in2 => \N__2678\,
            in3 => \N__2312\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNITMPMZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2309\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => \un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2300\,
            in3 => \N__2569\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_8_c_RNI3O5C_0_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2674\,
            lcout => \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_7_c_RNI1L4C_0_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2693\,
            lcout => \un5_visibley_cry_7_c_RNI1L4CZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_7_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__2427\,
            in1 => \N__3081\,
            in2 => \N__2333\,
            in3 => \N__2455\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4053\,
            ce => \N__2659\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__2360\,
            in1 => \N__2453\,
            in2 => \N__2429\,
            in3 => \N__3079\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4053\,
            ce => \N__2659\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__2426\,
            in1 => \N__3080\,
            in2 => \N__2351\,
            in3 => \N__2454\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4053\,
            ce => \N__2659\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3078\,
            in1 => \N__2428\,
            in2 => \N__2459\,
            in3 => \N__2483\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4053\,
            ce => \N__2659\,
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4146\,
            in2 => \N__2396\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => un21_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3041\,
            in2 => \_gnd_net_\,
            in3 => \N__2363\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => un21_beamy_cry_2,
            clk => \N__4052\,
            ce => \N__2666\,
            sr => \_gnd_net_\
        );

    \beamY_RNO_0_3_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2887\,
            in2 => \_gnd_net_\,
            in3 => \N__2354\,
            lcout => \beamY_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNO_0_4_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2857\,
            in2 => \_gnd_net_\,
            in3 => \N__2342\,
            lcout => \beamY_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_5_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2917\,
            in2 => \_gnd_net_\,
            in3 => \N__2339\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \N__4052\,
            ce => \N__2666\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2944\,
            in2 => \_gnd_net_\,
            in3 => \N__2336\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \N__4052\,
            ce => \N__2666\,
            sr => \_gnd_net_\
        );

    \beamY_RNO_0_7_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3117\,
            in2 => \_gnd_net_\,
            in3 => \N__2324\,
            lcout => \beamY_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_8_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2772\,
            in2 => \_gnd_net_\,
            in3 => \N__2321\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \N__4052\,
            ce => \N__2666\,
            sr => \_gnd_net_\
        );

    \beamY_RNO_0_9_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__2803\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2486\,
            lcout => \beamY_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3001\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2646\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIA525_0_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__2387\,
            in1 => \_gnd_net_\,
            in2 => \N__3152\,
            in3 => \N__3128\,
            lcout => un5_beamx_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNICPU5_1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3596\,
            in1 => \N__3233\,
            in2 => \N__3521\,
            in3 => \N__2968\,
            lcout => OPEN,
            ltout => \un3_beamx_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIKVE6_0_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3556\,
            in1 => \N__3419\,
            in2 => \N__2474\,
            in3 => \N__3000\,
            lcout => un3_beamx_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI5457_5_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__2471\,
            in1 => \N__3458\,
            in2 => \N__3638\,
            in3 => \N__3323\,
            lcout => \beamX_RNI5457Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIC725_9_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4141\,
            in1 => \N__2773\,
            in2 => \N__3047\,
            in3 => \N__2804\,
            lcout => un5_beamx_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__3082\,
            in1 => \N__2465\,
            in2 => \N__2422\,
            in3 => \N__2443\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4048\,
            ce => \N__2660\,
            sr => \_gnd_net_\
        );

    \beamY_0_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__2442\,
            in1 => \N__2409\,
            in2 => \N__2395\,
            in3 => \N__3083\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4048\,
            ce => \N__2660\,
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3005\,
            in2 => \N__2972\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3230\,
            in2 => \_gnd_net_\,
            in3 => \N__2510\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__4047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3551\,
            in2 => \_gnd_net_\,
            in3 => \N__2507\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__4047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2664\,
            in1 => \N__3592\,
            in2 => \_gnd_net_\,
            in3 => \N__2504\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__4047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3631\,
            in2 => \_gnd_net_\,
            in3 => \N__2501\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__4047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3410\,
            in2 => \_gnd_net_\,
            in3 => \N__2498\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__4047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3453\,
            in2 => \_gnd_net_\,
            in3 => \N__2495\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__4047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3365\,
            in2 => \_gnd_net_\,
            in3 => \N__2492\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__4047\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3343\,
            in2 => \_gnd_net_\,
            in3 => \N__2489\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__4046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2665\,
            in1 => \N__3506\,
            in2 => \_gnd_net_\,
            in3 => \N__2621\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2732\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2519\,
            in2 => \N__2547\,
            in3 => \N__2618\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5UR_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2540\,
            in2 => \N__2615\,
            in3 => \N__2606\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNID5URZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9K61_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2603\,
            in2 => \N__2548\,
            in3 => \N__2597\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIA9KZ0Z61\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNIVBNM1_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3275\,
            in1 => \N__2594\,
            in2 => \N__2588\,
            in3 => \N__2579\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2576\,
            in1 => \N__2568\,
            in2 => \N__2549\,
            in3 => \N__2525\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2522\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2710\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2731\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_2_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3046\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => un5_visibley_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_2_c_RNIN5VB_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2888\,
            in3 => \N__2741\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum\,
            ltout => OPEN,
            carryin => un5_visibley_cry_2,
            carryout => un5_visibley_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_3_c_RNIP80C_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2858\,
            in3 => \N__2738\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum\,
            ltout => OPEN,
            carryin => un5_visibley_cry_3,
            carryout => un5_visibley_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_4_c_RNIRB1C_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4297\,
            in2 => \N__2918\,
            in3 => \N__2735\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum\,
            ltout => OPEN,
            carryin => un5_visibley_cry_4,
            carryout => un5_visibley_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_5_c_RNITE2C_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4289\,
            in2 => \N__2945\,
            in3 => \N__2717\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum\,
            ltout => OPEN,
            carryin => un5_visibley_cry_5,
            carryout => un5_visibley_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_6_c_RNIVH3C_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4298\,
            in2 => \N__3120\,
            in3 => \N__2696\,
            lcout => \un1_beamY_if_generate_plus_mult1_un40_sum\,
            ltout => OPEN,
            carryin => un5_visibley_cry_6,
            carryout => un5_visibley_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_7_c_RNI1L4C_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4290\,
            in2 => \N__2774\,
            in3 => \N__2684\,
            lcout => \un5_visibley_cry_7_c_RNI1L4CZ0\,
            ltout => OPEN,
            carryin => un5_visibley_cry_7,
            carryout => un5_visibley_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_8_c_RNI3O5C_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2792\,
            in2 => \_gnd_net_\,
            in3 => \N__2681\,
            lcout => \un1_beamY_if_generate_plus_mult1_un33_sum_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__4299\,
            in1 => \N__3038\,
            in2 => \_gnd_net_\,
            in3 => \N__4177\,
            lcout => un5_visibley_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN4H2_5_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2942\,
            in2 => \_gnd_net_\,
            in3 => \N__2915\,
            lcout => un1_beamy_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_18_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3039\,
            in2 => \_gnd_net_\,
            in3 => \N__2884\,
            lcout => OPEN,
            ltout => \un4_beamylt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_14_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2943\,
            in1 => \N__2916\,
            in2 => \N__2894\,
            in3 => \N__2855\,
            lcout => OPEN,
            ltout => \un4_beamylt8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_5_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__2801\,
            in1 => \N__2771\,
            in2 => \N__2891\,
            in3 => \N__3118\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0H2_3_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2885\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2854\,
            lcout => un5_beamx_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_RNO_0_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__3119\,
            in1 => \N__3040\,
            in2 => \N__4151\,
            in3 => \N__2886\,
            lcout => OPEN,
            ltout => \un1_beamylto9_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__3167\,
            in1 => \N__3150\,
            in2 => \N__2861\,
            in3 => \N__2856\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITAH2_9_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2802\,
            in2 => \_gnd_net_\,
            in3 => \N__2770\,
            lcout => un8_beamy_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_7_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__3179\,
            in1 => \N__3634\,
            in2 => \N__3377\,
            in3 => \N__3595\,
            lcout => un18_beamylt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIQCL_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__2967\,
            in1 => \N__2999\,
            in2 => \N__3557\,
            in3 => \N__3232\,
            lcout => un18_beamylt4,
            ltout => \un18_beamylt4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_15_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101010101"
        )
    port map (
            in0 => \N__3418\,
            in1 => \N__3633\,
            in2 => \N__3173\,
            in3 => \N__3594\,
            lcout => OPEN,
            ltout => \un13_beamylt7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_6_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__3520\,
            in1 => \N__3322\,
            in2 => \N__3170\,
            in3 => \N__3457\,
            lcout => un13_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_13_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3163\,
            in1 => \N__3151\,
            in2 => \_gnd_net_\,
            in3 => \N__3127\,
            lcout => OPEN,
            ltout => \un8_beamylto9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_4_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000101"
        )
    port map (
            in0 => \N__3519\,
            in1 => \N__3072\,
            in2 => \N__3050\,
            in3 => \N__3042\,
            lcout => \Pixel_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2997\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => un5_visiblex_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__2998\,
            in1 => \N__2966\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_0,
            carryout => un5_visiblex_cry_1,
            clk => \N__4051\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3231\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => un5_visiblex_cry_1,
            carryout => un5_visiblex_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_9_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3544\,
            in2 => \N__4330\,
            in3 => \N__3203\,
            lcout => un1_visiblex_24,
            ltout => OPEN,
            carryin => un5_visiblex_cry_2,
            carryout => un5_visiblex_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3583\,
            in2 => \_gnd_net_\,
            in3 => \N__3200\,
            lcout => un1_visiblex_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_3,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3622\,
            in2 => \_gnd_net_\,
            in3 => \N__3197\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3400\,
            in2 => \N__4331\,
            in3 => \N__3194\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3447\,
            in2 => \_gnd_net_\,
            in3 => \N__3191\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3362\,
            in2 => \N__4332\,
            in3 => \N__3188\,
            lcout => \un5_visiblex_cry_7_c_RNIVZ0Z952\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3338\,
            in2 => \_gnd_net_\,
            in3 => \N__3185\,
            lcout => un1_visiblex_if_generate_plus_mult1_un40_sum_c5,
            ltout => \un1_visiblex_if_generate_plus_mult1_un40_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3182\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un40_sum_c5_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_RNO_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3632\,
            in1 => \N__3593\,
            in2 => \N__3411\,
            in3 => \N__3552\,
            lcout => OPEN,
            ltout => \un1_beamxlt10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__3507\,
            in1 => \N__3321\,
            in2 => \N__3485\,
            in3 => \N__3449\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_16_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3364\,
            in1 => \N__3448\,
            in2 => \N__3344\,
            in3 => \N__3401\,
            lcout => un18_beamylto9_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIR4B_9_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3339\,
            lcout => un1_beamx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3833\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3276\,
            in2 => \N__3302\,
            in3 => \N__3293\,
            lcout => \un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3290\,
            in2 => \N__3281\,
            in3 => \N__3284\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8IL1_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3280\,
            in2 => \N__3260\,
            in3 => \N__3251\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNIT8ILZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQ5N04_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3692\,
            in1 => \N__3248\,
            in2 => \N__3242\,
            in3 => \N__3725\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3722\,
            in2 => \_gnd_net_\,
            in3 => \N__3716\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02\,
            ltout => \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMDZ0Z02_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNIVMD02_0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3713\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3946\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFR2_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3693\,
            in2 => \N__3818\,
            in3 => \N__3710\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIATFRZ0Z2\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6B3_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3707\,
            in2 => \N__3698\,
            in3 => \N__3701\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIRJ6BZ0Z3\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3R3_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3697\,
            in2 => \N__3677\,
            in3 => \N__3668\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIAJ3RZ0Z3\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIHBHM8_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3791\,
            in1 => \N__3665\,
            in2 => \N__3659\,
            in3 => \N__3650\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3647\,
            in2 => \_gnd_net_\,
            in3 => \N__3641\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4\,
            ltout => \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKGZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNIOPKG4_0_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3836\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3832\,
            lcout => \un1_beamY_if_generate_plus_mult1_un54_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3737\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3O4_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3792\,
            in2 => \N__3935\,
            in3 => \N__3809\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNI8V3OZ0Z4\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFE7_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3806\,
            in2 => \N__3797\,
            in3 => \N__3800\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNI4PFEZ0Z7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7U7_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3796\,
            in2 => \N__3776\,
            in3 => \N__3767\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNIMH7UZ0Z7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNIS657H_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3888\,
            in1 => \N__3764\,
            in2 => \N__3758\,
            in3 => \N__3749\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_axb_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVO8_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3746\,
            in2 => \_gnd_net_\,
            in3 => \N__3740\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMJVOZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3947\,
            lcout => \un1_beamY_if_generate_plus_mult1_un61_sum_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_17_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4173\,
            in2 => \_gnd_net_\,
            in3 => \N__4145\,
            lcout => \G_6_i_a4_0_0\,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFP59_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3926\,
            in2 => \N__3889\,
            in3 => \N__3920\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNIBFPZ0Z59\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_2\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPD_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3884\,
            in2 => \N__3917\,
            in3 => \N__3908\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNIUTLPDZ0\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_3\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_12_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3905\,
            in2 => \N__3890\,
            in3 => \N__3899\,
            lcout => \Pixel_1_RNOZ0Z_12\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_4\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3896\,
            in2 => \N__3863\,
            in3 => \N__3880\,
            lcout => \un1_beamY_if_generate_plus_mult1_un68_sum_i_7\,
            ltout => OPEN,
            carryin => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_5\,
            carryout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFH_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3854\,
            in2 => \_gnd_net_\,
            in3 => \N__3848\,
            lcout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0\,
            ltout => \un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNIVNQFHZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_11_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3845\,
            in1 => \N__4202\,
            in2 => \N__3839\,
            in3 => \N__4190\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_10_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4201\,
            in1 => \N__4189\,
            in2 => \N__4178\,
            in3 => \N__4157\,
            lcout => OPEN,
            ltout => \N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110100"
        )
    port map (
            in0 => \N__4150\,
            in1 => \N__4100\,
            in2 => \N__4094\,
            in3 => \N__4091\,
            lcout => OPEN,
            ltout => \un15_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000100"
        )
    port map (
            in0 => \N__3956\,
            in1 => \N__3986\,
            in2 => \N__4085\,
            in3 => \N__3965\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4019\,
            in1 => \N__4013\,
            in2 => \N__4007\,
            in3 => \N__3995\,
            lcout => \Pixel_0_sqmuxa_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4530\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_2_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100010100010"
        )
    port map (
            in0 => \N__4418\,
            in1 => \N__4450\,
            in2 => \N__3980\,
            in3 => \N__4634\,
            lcout => un14lt10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_1_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100111001100"
        )
    port map (
            in0 => \N__4417\,
            in1 => \N__4406\,
            in2 => \N__4451\,
            in3 => \N__4633\,
            lcout => un1_visiblex_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4381\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUK_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4502\,
            in2 => \N__4460\,
            in3 => \N__4397\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNIGUUKZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBM831_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4492\,
            in2 => \N__4358\,
            in3 => \N__4394\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIBMZ0Z831\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISON62_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4691\,
            in1 => \N__4478\,
            in2 => \N__4214\,
            in3 => \N__4391\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4493\,
            in1 => \N__4541\,
            in2 => \N__4517\,
            in3 => \N__4388\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUCZ0Z31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIFUC31_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4385\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4382\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4471\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDG_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4367\,
            in2 => \_gnd_net_\,
            in3 => \N__4349\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNIPVDGZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FG_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4346\,
            in2 => \N__4337\,
            in3 => \N__4205\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQ1FGZ0\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4537\,
            in2 => \_gnd_net_\,
            in3 => \N__4508\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4505\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4496\,
            in3 => \_gnd_net_\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4481\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4472\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un5_visiblex_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4446\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2G5_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4645\,
            in2 => \N__4625\,
            in3 => \N__4409\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_RNII2GZ0Z5\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_8_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4592\,
            in2 => \N__4559\,
            in3 => \N__4400\,
            lcout => \Pixel_1_RNOZ0Z_8\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4646\,
            in2 => \N__4583\,
            in3 => \N__4554\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PB_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4571\,
            in2 => \_gnd_net_\,
            in3 => \N__4637\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_RNIC20PBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4616\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4615\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90R03_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4711\,
            in2 => \N__4655\,
            in3 => \N__4586\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNI90RZ0Z03\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80F4_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4727\,
            in2 => \N__4778\,
            in3 => \N__4574\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIF80FZ0Z4\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6_c_RNIGQELB_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4558\,
            in1 => \N__4712\,
            in2 => \N__4757\,
            in3 => \N__4565\,
            lcout => un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJ6_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4745\,
            in2 => \_gnd_net_\,
            in3 => \N__4562\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNICMHJZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4670\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_6_0_\,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7G1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4793\,
            in2 => \N__4787\,
            in3 => \N__4769\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI0A7GZ0Z1\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIK3332_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4690\,
            in2 => \N__4766\,
            in3 => \N__4748\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKZ0Z3332\,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNIEN766_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4726\,
            in1 => \N__4676\,
            in2 => \N__4703\,
            in3 => \N__4739\,
            lcout => un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4736\,
            in2 => \_gnd_net_\,
            in3 => \N__4730\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2\,
            ltout => \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HHZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJ3HH2_0_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4715\,
            in3 => \_gnd_net_\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKL62_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4702\,
            in2 => \_gnd_net_\,
            in3 => \N__4689\,
            lcout => \un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIQKLZ0Z62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4669\,
            lcout => un1_visiblex_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
