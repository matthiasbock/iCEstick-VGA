-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 23 2015 22:12:10

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__16788\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16463\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16325\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16268\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16135\ : std_logic;
signal \N__16132\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16091\ : std_logic;
signal \N__16088\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16052\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15781\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15707\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15347\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14403\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14111\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13760\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13727\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13718\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13694\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13241\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7275\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_4_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2_cascade_\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRUZ0Z85\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDCZ0Z3\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PUZ0Z3\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJZ0Z4\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8AZ0Z6\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RHZ0Z9\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74AZ0\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal \chary_if_generate_plus_mult1_un47_sum_axb4_cascade_\ : std_logic;
signal \beamY_RNIKM9GCZ0Z_9_cascade_\ : std_logic;
signal \beamY_RNIM5433Z0Z_8\ : std_logic;
signal \beamY_RNI93821Z0Z_9_cascade_\ : std_logic;
signal \beamY_RNIM5433_0Z0Z_8\ : std_logic;
signal \beamY_RNIIR4K3_0Z0Z_7\ : std_logic;
signal \beamY_RNIIR4K3_0Z0Z_7_cascade_\ : std_logic;
signal \beamY_RNIKM9GC_0Z0Z_9\ : std_logic;
signal \chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_\ : std_logic;
signal \beamY_RNI9DSP2_0Z0Z_8\ : std_logic;
signal \beamY_RNI41384Z0Z_7_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un54_sum_ac0_5_1_cascade_\ : std_logic;
signal \un8_beamylt9_0_cascade_\ : std_logic;
signal \beamY_RNIP8FF1_1Z0Z_7\ : std_logic;
signal \beamY_RNI93821Z0Z_9\ : std_logic;
signal \beamY_RNIBV5E51Z0Z_8_cascade_\ : std_logic;
signal \beamY_RNIBV5E51_0Z0Z_8\ : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_axbxc5_2 : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_c5 : std_logic;
signal \beamY_RNIVADQVZ0Z_8_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_ac0_5 : std_logic;
signal \beamY_RNIV5SUC3_0Z0Z_9_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb4_0_1 : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_axb4_0_cascade_\ : std_logic;
signal \beamY_RNIVADQVZ0Z_8\ : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_c4 : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_axb4 : std_logic;
signal \beamY_RNIV5SUC3Z0Z_9\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_0 : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_axb4_0_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_axb4_i_cascade_\ : std_logic;
signal g1_0_2 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axb4_0 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axb4_i_0 : std_logic;
signal g1_1 : std_logic;
signal \g2_0_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_axb4_i_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__g0Z0Z_2\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb4_0 : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_c4_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb3_0 : std_logic;
signal \beamY_RNISDTA58Z0Z_5_cascade_\ : std_logic;
signal \beamY_RNIJ0797KZ0Z_4\ : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal \beamY_RNI2B511_0Z0Z_9\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \beamY_RNIUUEM_0Z0Z_8\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVLZ0Z21\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1NZ0Z21\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal \bfn_2_4_0_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6UZ0\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVHZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEAZ0Z1\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8UZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HAZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_axb3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NEZ0\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATKZ0\ : std_logic;
signal \beamY_i_2_cascade_\ : std_logic;
signal \beamY_fast_RNIT5UFZ0Z_4_cascade_\ : std_logic;
signal un5_visibley_ac0_7 : std_logic;
signal \un5_visibley_ac0_7_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux : std_logic;
signal \beamY_fastZ0Z_7\ : std_logic;
signal \beamY_fastZ0Z_6\ : std_logic;
signal \beamY_fastZ0Z_5\ : std_logic;
signal \un5_visibley_ac0_11_0_1_cascade_\ : std_logic;
signal \beamY_fastZ0Z_4\ : std_logic;
signal \beamY_fastZ0Z_8\ : std_logic;
signal un5_visibley_c7 : std_logic;
signal \beamY_fastZ0Z_3\ : std_logic;
signal \un5_visibley_c2_cascade_\ : std_logic;
signal \beamY_fastZ0Z_2\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \un21_beamy_cry_1_c_RNIALZ0Z73\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal \un21_beamy_cry_2_c_RNICOZ0Z83\ : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal \un21_beamy_cry_3_c_RNIERZ0Z93\ : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal \un21_beamy_cry_4_c_RNIGUAZ0Z3\ : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal \un21_beamy_cry_5_c_RNII1CZ0Z3\ : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal \un21_beamy_cry_6_c_RNIK4DZ0Z3\ : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal \un21_beamy_cry_7_c_RNIM7EZ0Z3\ : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal \bfn_2_13_0_\ : std_logic;
signal \if_generate_plus_mult1_un61_sum_axbxc5_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_ac0_7_dZ0_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_c5_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un61_sum_axb4_i : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_6\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_ac0_7_0Z0Z_1\ : std_logic;
signal \row_1_if_i4_mux_i_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\ : std_logic;
signal row_1_if_i4_mux_i : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_ac0_7_0Z0Z_1_cascade_\ : std_logic;
signal \row_1_if_N_6\ : std_logic;
signal \if_generate_plus_mult1_un75_sum_axbxc3_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0\ : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0\ : std_logic;
signal if_generate_plus_mult1_un75_sum_axbxc3 : std_logic;
signal row_1_if_generate_plus_mult1_un75_sum_c5 : std_logic;
signal \if_generate_plus_mult1_un82_sum_axb4_x1_cascade_\ : std_logic;
signal if_generate_plus_mult1_un82_sum_axb4_x0 : std_logic;
signal \beamY_RNIP8FF1_0Z0Z_7\ : std_logic;
signal \un114_pixel_6_1_5__un5_beamxZ0Z_3_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__un5_beamxZ0Z_5_cascade_\ : std_logic;
signal \beamY_RNIP8FF1Z0Z_7_cascade_\ : std_logic;
signal un5_visibley_c6 : std_logic;
signal chary_if_generate_plus_mult1_un40_sum_c4 : std_logic;
signal un5_visibley_c5 : std_logic;
signal \beamY_RNIP8FF1_2Z0Z_7\ : std_logic;
signal \un4_beamylt6_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_axbxc5_1 : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_c5 : std_logic;
signal \beamY_RNIB6AOI5_0Z0Z_5_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_7_d : std_logic;
signal un5_visibley_c2 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum : std_logic;
signal g2_1 : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_c5_0_cascade_\ : std_logic;
signal \chary_if_generate_plus_mult1_un1_sum_axbxc3_1_1_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_axb3 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axbxc5_0 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c5_0_0 : std_logic;
signal \un114_pixel_6_1_5__g0_17Z0Z_1_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un75_sum_0_5 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb4_i : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_c4 : std_logic;
signal g1_0_3 : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal row_1_if_generate_plus_mult1_un82_sum_axb4_i : std_logic;
signal \un114_pixel_6_1_5__un8_beamylto9Z0Z_0\ : std_logic;
signal un8_beamylt9_0 : std_logic;
signal \un114_pixel_6_1_5__un1_beamylto9Z0Z_0_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__un1_beamylto9_3_cascade_\ : std_logic;
signal \VSync_c\ : std_logic;
signal un8_beamy_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un61_sum_c5 : std_logic;
signal \row_1_if_generate_plus_mult1_un82_sum_axbxc5_3Z0Z_1_cascade_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum : std_logic;
signal un4_beamylt8_0 : std_logic;
signal \un114_pixel_6_1_5__g0_1Z0Z_4_cascade_\ : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal \un114_pixel_6_1_5__g0_0Z0Z_4\ : std_logic;
signal \un114_pixel_6_1_5__g0_0Z0Z_3_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__g2_0Z0Z_0_cascade_\ : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \un114_pixel_6_1_5__g0_0_1Z0Z_1\ : std_logic;
signal g1 : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cascade_\ : std_logic;
signal m511_0_x2_1_2 : std_logic;
signal \G_7_0_m2_1_1_1_cascade_\ : std_logic;
signal \G_7_0_m2_1_1_cascade_\ : std_logic;
signal \G_7_0_m2_1_0\ : std_logic;
signal chary_if_generate_plus_mult1_un75_sum_c5 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c4 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_c5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axbxc5_1 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_ac0_5 : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_\ : std_logic;
signal \beamY_RNIL0E2QG2Z0Z_3\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal un5_visiblex_cry_0 : std_logic;
signal un5_visiblex_cry_1 : std_logic;
signal un5_visiblex_cry_2 : std_logic;
signal un5_visiblex_cry_3 : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axbxc5 : std_logic;
signal if_generate_plus_mult1_un61_sum_axbxc5 : std_logic;
signal \un114_pixel_6_1_5__un3_beamxZ0Z_5_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__un3_beamxZ0Z_7\ : std_logic;
signal \un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1Z0Z_1\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0\ : std_logic;
signal un4_beamy_0 : std_logic;
signal \un13_beamylt10_0_cascade_\ : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un18_beamylt5_0 : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal \un18_beamylt5_0_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__un15_beamyZ0Z_0\ : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal \un114_pixel_6_1_5__un18_beamylto9Z0Z_2\ : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal \un114_pixel_6_1_5__un13_beamylto2Z0Z_0\ : std_logic;
signal \un114_pixel_6_1_5__un15_beamyZ0Z_1\ : std_logic;
signal un4_beamy_0_0 : std_logic;
signal \un114_pixel_6_1_5__g3_0_0_0\ : std_logic;
signal un13_beamylt10_0 : std_logic;
signal un1_beamx_2 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal un1_beamxlt10_0 : std_logic;
signal \HSync_c\ : std_logic;
signal \un114_pixel_6_1_5__un4_rowZ0Z_5\ : std_logic;
signal row_1_if_generate_plus_mult1_un68_sum_c5 : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\ : std_logic;
signal if_generate_plus_mult1_un75_sum_axbxc5 : std_logic;
signal \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_3\ : std_logic;
signal \un114_pixel_6_1_5__un4_rowZ0Z_7_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__un4_rowZ0Z_1\ : std_logic;
signal \beamY_i_2\ : std_logic;
signal \un114_pixel_6_1_5__chessboardpixel_un200_pixellto4Z0Z_1\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4OZ0\ : std_logic;
signal \chessboardpixel_un200_pixellt10_cascade_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c5_0 : std_logic;
signal \chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_cascade_\ : std_logic;
signal g1_0_1 : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axb4_i : std_logic;
signal g2 : std_logic;
signal m511_0_o2_1 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axbxc5_0 : std_logic;
signal \N_80_i\ : std_logic;
signal un3_beamx_0 : std_logic;
signal un5_beamx_0 : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_0 : std_logic;
signal \beamY_RNIJH2N2PZ0Z_3\ : std_logic;
signal \bfn_7_3_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_2 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_4 : std_logic;
signal \column_1_if_generate_plus_mult1_un47_sum1_5_cascade_\ : std_logic;
signal un5_visiblex_i_0_25 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_axb_3_i : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_4 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_3 : std_logic;
signal \if_generate_plus_mult1_un47_sum_m_5_cascade_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_\ : std_logic;
signal \N_11_0_i\ : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3 : std_logic;
signal chary_if_generate_plus_mult1_un33_sum_axb3 : std_logic;
signal \un114_pixel_6_1_5__un4_rowZ0Z_2\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal if_generate_plus_mult1_un47_sum_m_1 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un47_sum_m_5 : std_logic;
signal if_generate_plus_mult1_un47_sum_m_2 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_4_l_fx : std_logic;
signal \N_571_i\ : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \if_generate_plus_mult1_un54_sum_s_5_cascade_\ : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un54_sum_s_5 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \N_562_i\ : std_logic;
signal chessboardpixel_un174_pixel_0_1 : std_logic;
signal chessboardpixel_un200_pixel_0_1 : std_logic;
signal \un114_pixel_6_1_5__un4_row_7Z0Z_1\ : std_logic;
signal \N_357_0\ : std_logic;
signal \N_18_0_cascade_\ : std_logic;
signal \N_7_0_cascade_\ : std_logic;
signal font_un28_pixel_0_0_29 : std_logic;
signal \un114_pixel_6_1_5__un116_pixel_3_1_0_0_7_cascade_\ : std_logic;
signal \N_14_0\ : std_logic;
signal \column_0111_0_cascade_\ : std_logic;
signal \beamY_RNI05CI5A3_0Z0Z_0_cascade_\ : std_logic;
signal \beamY_RNIBABJS01Z0Z_1_cascade_\ : std_logic;
signal \N_21_0_cascade_\ : std_logic;
signal \N_22_0\ : std_logic;
signal column_0111_0 : std_logic;
signal \un116_pixel_3_bmZ0Z_6_cascade_\ : std_logic;
signal \beamY_RNISJITRQ2Z0Z_1_cascade_\ : std_logic;
signal \N_12_0\ : std_logic;
signal \N_248_0_cascade_\ : std_logic;
signal un116_pixel_3_ns_1_0_6 : std_logic;
signal \N_25_mux\ : std_logic;
signal \un114_pixel_3_i_a3_7_cascade_\ : std_logic;
signal column_0001_0 : std_logic;
signal \un116_pixel_3_ns_1_2_cascade_\ : std_logic;
signal \beamY_RNIDVSK5A3Z0Z_1\ : std_logic;
signal \N_13_0\ : std_logic;
signal \un114_pixel_0_1__N_6_mux_0\ : std_logic;
signal \un116_pixel_1_amZ0Z_1_cascade_\ : std_logic;
signal \un116_pixel_4_bmZ0Z_1\ : std_logic;
signal \un116_pixel_4_amZ0Z_1_cascade_\ : std_logic;
signal un116_pixel_3_ns_1_1 : std_logic;
signal \beamY_RNIHIRVUS1Z0Z_1\ : std_logic;
signal \un116_pixel_1_bmZ0Z_1\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_2 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_2 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_4 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_4 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_cry_3_ma : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx : std_logic;
signal \N_200_0_i\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_s_2_sf : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_1 : std_logic;
signal \un5_visiblex_cry_8_c_RNI1D62Z0Z_2\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_4 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx : std_logic;
signal un5_visiblex_i_25 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_5 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_5 : std_logic;
signal \un114_pixel_6_1_5__un4_rowZ0Z_0\ : std_logic;
signal \un116_pixel_5_amZ0Z_6_cascade_\ : std_logic;
signal \un116_pixel_5_bmZ0Z_6\ : std_logic;
signal un15_beamy : std_logic;
signal \un114_pixel_6_1_5__g0Z0Z_0\ : std_logic;
signal \un114_pixel_6_1_5__font_un126_pixel_mZ0Z_1_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__font_un126_pixel_m_4_1_0\ : std_logic;
signal \un114_pixel_6_1_5__g0_2Z0Z_0_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__font_un126_pixel_m_4_1_1_0\ : std_logic;
signal \un114_pixel_6_1_5__g0_1_0\ : std_logic;
signal \un114_pixel_6_1_5__g1Z0Z_0_cascade_\ : std_logic;
signal un4_row : std_logic;
signal \beamY_RNIPG1SS93Z0Z_2\ : std_logic;
signal \N_23_0\ : std_logic;
signal \N_15_0\ : std_logic;
signal \N_342_0_0\ : std_logic;
signal \N_1045_0_cascade_\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_iZ0\ : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal un5_rowlto3_i : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \Pixel_3_sqmuxa\ : std_logic;
signal \un114_pixel_6_1_5__font_un126_pixel_m_4\ : std_logic;
signal un1_beamy_0_0 : std_logic;
signal \Pixel_1_r_sn\ : std_logic;
signal \Pixel_1_r_rn_0_cascade_\ : std_logic;
signal \N_396\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal \m6Z0Z_1\ : std_logic;
signal \G_7_0_m2_1\ : std_logic;
signal \beamX_RNI1M3Q1V2Z0Z_0_cascade_\ : std_logic;
signal \N_1039_0_0\ : std_logic;
signal \font_un3_pixel_29_cascade_\ : std_logic;
signal \G_7_0_m4_2_1_1_cascade_\ : std_logic;
signal \G_7_0_m4_2_1\ : std_logic;
signal \beamY_RNINIKJ5A3Z0Z_1\ : std_logic;
signal \beamY_RNI7OTDJ61Z0Z_1_cascade_\ : std_logic;
signal \beamY_RNIJDHE4C2Z0Z_1\ : std_logic;
signal \font_un126_pixel_6_am_cascade_\ : std_logic;
signal font_un126_pixel_2_am : std_logic;
signal \beamX_RNIQ6MATS2Z0Z_0\ : std_logic;
signal \un114_pixel_7_1_7__N_11_i_1\ : std_logic;
signal \N_37_cascade_\ : std_logic;
signal \beamY_RNI05CI5A3_1Z0Z_0_cascade_\ : std_logic;
signal \beamY_RNI05CI5A3Z0Z_0\ : std_logic;
signal \beamY_RNII25UDD3_1Z0Z_0\ : std_logic;
signal \un116_pixel_7_ns_1_4_cascade_\ : std_logic;
signal \beamY_RNIFHEQCT1Z0Z_0\ : std_logic;
signal \beamY_RNIA4V0NM1Z0Z_0_cascade_\ : std_logic;
signal \beamY_RNII25UDD3_0Z0Z_0\ : std_logic;
signal \un116_pixel_7_ns_1_6_cascade_\ : std_logic;
signal font_un3_pixel_29 : std_logic;
signal \beamY_RNIBHJ7AMZ0Z_0\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_iZ0\ : std_logic;
signal \G_340\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_2 : std_logic;
signal \G_341\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_4 : std_logic;
signal \un5_rowlto0_cascade_\ : std_logic;
signal \beamY_RNIJ720T72Z0Z_0\ : std_logic;
signal un116_pixel_5_ns_1_2 : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_iZ0\ : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_2_s : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un116_pixel_2_ns_1_2 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_3_s : std_logic;
signal if_generate_plus_mult1_un75_sum_axb_4_l_fx : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0\ : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum : std_logic;
signal \N_520\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal un5_visiblex_i_24 : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal \CO3_0\ : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0_cascade_\ : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\ : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_\ : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4 : std_logic;
signal \un114_pixel_6_1_5__g2_0_1\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPBZ0Z3\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__font_un126_pixel_m_1Z0Z_1\ : std_logic;
signal charx_if_generate_plus_mult1_un1_sum_axb1 : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\ : std_logic;
signal \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__font_un126_pixel_m_1_1Z0Z_1\ : std_logic;
signal \m15_cascade_\ : std_logic;
signal \un114_pixel_0_1__N_6_mux\ : std_logic;
signal \beamY_RNI4NRC8D1Z0Z_0_cascade_\ : std_logic;
signal \beamY_RNII25UDD3Z0Z_0\ : std_logic;
signal \N_14\ : std_logic;
signal \un116_pixel_2_ns_1_6_cascade_\ : std_logic;
signal \beamY_RNIH01F2SZ0Z_0\ : std_logic;
signal \un116_pixel_2_ns_1Z0Z_5\ : std_logic;
signal \N_276_0_cascade_\ : std_logic;
signal \beamY_RNII25UDD3_3Z0Z_0\ : std_logic;
signal m7 : std_logic;
signal \m7_cascade_\ : std_logic;
signal \N_302_i_0\ : std_logic;
signal \beamY_RNITQPUS72Z0Z_0_cascade_\ : std_logic;
signal un116_pixel_3_1_0 : std_logic;
signal \beamY_RNI6B7UAL1Z0Z_1\ : std_logic;
signal m31 : std_logic;
signal \un116_pixel_4_1Z0Z_0\ : std_logic;
signal m38 : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal \m38_cascade_\ : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal \un116_pixel_6_1_1_cascade_\ : std_logic;
signal \N_17\ : std_logic;
signal \N_321\ : std_logic;
signal \un116_pixel_2_bmZ0Z_1\ : std_logic;
signal un5_rowlto2_i : std_logic;
signal un5_rowlto2 : std_logic;
signal un5_rowlto0 : std_logic;
signal un5_rowlto1 : std_logic;
signal un5_rowlto3 : std_logic;
signal \un116_pixel_2_amZ0Z_1\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\ : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\ : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\ : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal chessboardpixel_un152_pixel_24 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal charx_i_24 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3Z0Z_0\ : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf : std_logic;
signal charx_i_23 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \PixelDebug_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    Pixel <= \Pixel_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    HSyncDebug <= \HSyncDebug_wire\;
    PixelDebug <= \PixelDebug_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__6839\,
            RESETB => \N__14250\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16788\,
            DIN => \N__16787\,
            DOUT => \N__16786\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16788\,
            PADOUT => \N__16787\,
            PADIN => \N__16786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9202\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16779\,
            DIN => \N__16778\,
            DOUT => \N__16777\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16779\,
            PADOUT => \N__16778\,
            PADIN => \N__16777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11098\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16770\,
            DIN => \N__16769\,
            DOUT => \N__16768\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16770\,
            PADOUT => \N__16769\,
            PADIN => \N__16768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13178\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16761\,
            DIN => \N__16760\,
            DOUT => \N__16759\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16761\,
            PADOUT => \N__16760\,
            PADIN => \N__16759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9209\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16752\,
            DIN => \N__16751\,
            DOUT => \N__16750\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__16752\,
            PADOUT => \N__16751\,
            PADIN => \N__16750\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16743\,
            DIN => \N__16742\,
            DOUT => \N__16741\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16743\,
            PADOUT => \N__16742\,
            PADIN => \N__16741\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11102\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16734\,
            DIN => \N__16733\,
            DOUT => \N__16732\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16734\,
            PADOUT => \N__16733\,
            PADIN => \N__16732\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13177\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3889\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16712\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__16712\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__16709\,
            I => \N__16705\
        );

    \I__3886\ : InMux
    port map (
            O => \N__16708\,
            I => \N__16701\
        );

    \I__3885\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16696\
        );

    \I__3884\ : InMux
    port map (
            O => \N__16704\,
            I => \N__16696\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__16701\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__16696\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__16691\,
            I => \N__16687\
        );

    \I__3880\ : CascadeMux
    port map (
            O => \N__16690\,
            I => \N__16684\
        );

    \I__3879\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16679\
        );

    \I__3878\ : InMux
    port map (
            O => \N__16684\,
            I => \N__16679\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__16679\,
            I => charx_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3875\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__16670\,
            I => charx_if_generate_plus_mult1_un75_sum_axb_5
        );

    \I__3873\ : InMux
    port map (
            O => \N__16667\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__3871\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16658\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__16658\,
            I => \N__16655\
        );

    \I__3869\ : Odrv4
    port map (
            O => \N__16655\,
            I => charx_i_24
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__16652\,
            I => \N__16649\
        );

    \I__3867\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16646\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__16646\,
            I => \N__16643\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__16643\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3Z0Z_0\
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__16640\,
            I => \N__16636\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__16639\,
            I => \N__16632\
        );

    \I__3862\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16625\
        );

    \I__3861\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16625\
        );

    \I__3860\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16625\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__16625\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\
        );

    \I__3858\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16618\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__16621\,
            I => \N__16615\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__16618\,
            I => \N__16612\
        );

    \I__3855\ : InMux
    port map (
            O => \N__16615\,
            I => \N__16609\
        );

    \I__3854\ : Span4Mux_h
    port map (
            O => \N__16612\,
            I => \N__16606\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__16609\,
            I => \N__16603\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__16606\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__3851\ : Odrv4
    port map (
            O => \N__16603\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__16598\,
            I => \N__16595\
        );

    \I__3849\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16592\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__16592\,
            I => \N__16589\
        );

    \I__3847\ : Span4Mux_h
    port map (
            O => \N__16589\,
            I => \N__16586\
        );

    \I__3846\ : Odrv4
    port map (
            O => \N__16586\,
            I => charx_i_23
        );

    \I__3845\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16574\
        );

    \I__3844\ : InMux
    port map (
            O => \N__16582\,
            I => \N__16563\
        );

    \I__3843\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16563\
        );

    \I__3842\ : InMux
    port map (
            O => \N__16580\,
            I => \N__16563\
        );

    \I__3841\ : InMux
    port map (
            O => \N__16579\,
            I => \N__16563\
        );

    \I__3840\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16563\
        );

    \I__3839\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16559\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__16574\,
            I => \N__16556\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__16563\,
            I => \N__16553\
        );

    \I__3836\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16550\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__16559\,
            I => \N__16547\
        );

    \I__3834\ : Span4Mux_v
    port map (
            O => \N__16556\,
            I => \N__16544\
        );

    \I__3833\ : Span4Mux_h
    port map (
            O => \N__16553\,
            I => \N__16539\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__16550\,
            I => \N__16539\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__16547\,
            I => \N__16536\
        );

    \I__3830\ : Span4Mux_v
    port map (
            O => \N__16544\,
            I => \N__16531\
        );

    \I__3829\ : Span4Mux_v
    port map (
            O => \N__16539\,
            I => \N__16531\
        );

    \I__3828\ : Span4Mux_v
    port map (
            O => \N__16536\,
            I => \N__16528\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__16531\,
            I => \N__16525\
        );

    \I__3826\ : Odrv4
    port map (
            O => \N__16528\,
            I => charx_if_generate_plus_mult1_un75_sum
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__16525\,
            I => charx_if_generate_plus_mult1_un75_sum
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__16520\,
            I => \N__16517\
        );

    \I__3823\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16502\
        );

    \I__3822\ : InMux
    port map (
            O => \N__16516\,
            I => \N__16502\
        );

    \I__3821\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16502\
        );

    \I__3820\ : InMux
    port map (
            O => \N__16514\,
            I => \N__16502\
        );

    \I__3819\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16502\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__16502\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\
        );

    \I__3817\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16496\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__16496\,
            I => \N__16492\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__16495\,
            I => \N__16487\
        );

    \I__3814\ : Span4Mux_h
    port map (
            O => \N__16492\,
            I => \N__16482\
        );

    \I__3813\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16471\
        );

    \I__3812\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16471\
        );

    \I__3811\ : InMux
    port map (
            O => \N__16487\,
            I => \N__16471\
        );

    \I__3810\ : InMux
    port map (
            O => \N__16486\,
            I => \N__16471\
        );

    \I__3809\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16471\
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__16482\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__16471\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\
        );

    \I__3806\ : CascadeMux
    port map (
            O => \N__16466\,
            I => \N__16463\
        );

    \I__3805\ : InMux
    port map (
            O => \N__16463\,
            I => \N__16460\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__16460\,
            I => \N__16457\
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__16457\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\
        );

    \I__3802\ : InMux
    port map (
            O => \N__16454\,
            I => \N__16451\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__16451\,
            I => \N__16448\
        );

    \I__3800\ : Span4Mux_v
    port map (
            O => \N__16448\,
            I => \N__16443\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__16447\,
            I => \N__16440\
        );

    \I__3798\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16436\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__16443\,
            I => \N__16433\
        );

    \I__3796\ : InMux
    port map (
            O => \N__16440\,
            I => \N__16430\
        );

    \I__3795\ : InMux
    port map (
            O => \N__16439\,
            I => \N__16427\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__16436\,
            I => \N__16424\
        );

    \I__3793\ : Sp12to4
    port map (
            O => \N__16433\,
            I => \N__16419\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__16430\,
            I => \N__16419\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__16427\,
            I => \N__16416\
        );

    \I__3790\ : Span4Mux_h
    port map (
            O => \N__16424\,
            I => \N__16413\
        );

    \I__3789\ : Span12Mux_s6_h
    port map (
            O => \N__16419\,
            I => \N__16410\
        );

    \I__3788\ : Odrv12
    port map (
            O => \N__16416\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__3787\ : Odrv4
    port map (
            O => \N__16413\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__3786\ : Odrv12
    port map (
            O => \N__16410\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__3785\ : InMux
    port map (
            O => \N__16403\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__3784\ : InMux
    port map (
            O => \N__16400\,
            I => \N__16396\
        );

    \I__3783\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16393\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__16396\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__16393\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__16388\,
            I => \N__16385\
        );

    \I__3779\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16382\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__16382\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7\
        );

    \I__3777\ : InMux
    port map (
            O => \N__16379\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__3776\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16373\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__16373\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__16370\,
            I => \N__16366\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__16369\,
            I => \N__16363\
        );

    \I__3772\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16358\
        );

    \I__3771\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16358\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__16358\,
            I => charx_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__3769\ : InMux
    port map (
            O => \N__16355\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__3768\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16349\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__16349\,
            I => charx_if_generate_plus_mult1_un68_sum_axb_5
        );

    \I__3766\ : InMux
    port map (
            O => \N__16346\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__3765\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16340\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__16340\,
            I => \N__16336\
        );

    \I__3763\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16333\
        );

    \I__3762\ : Span4Mux_v
    port map (
            O => \N__16336\,
            I => \N__16328\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__16333\,
            I => \N__16328\
        );

    \I__3760\ : Span4Mux_h
    port map (
            O => \N__16328\,
            I => \N__16322\
        );

    \I__3759\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16319\
        );

    \I__3758\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16316\
        );

    \I__3757\ : CascadeMux
    port map (
            O => \N__16325\,
            I => \N__16313\
        );

    \I__3756\ : Sp12to4
    port map (
            O => \N__16322\,
            I => \N__16306\
        );

    \I__3755\ : LocalMux
    port map (
            O => \N__16319\,
            I => \N__16306\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__16316\,
            I => \N__16306\
        );

    \I__3753\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16303\
        );

    \I__3752\ : Span12Mux_s11_v
    port map (
            O => \N__16306\,
            I => \N__16300\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__16303\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__3750\ : Odrv12
    port map (
            O => \N__16300\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__3749\ : InMux
    port map (
            O => \N__16295\,
            I => \N__16292\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__16292\,
            I => charx_if_generate_plus_mult1_un61_sum_i
        );

    \I__3747\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16286\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__16286\,
            I => \N__16283\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__16283\,
            I => charx_if_generate_plus_mult1_un68_sum_i
        );

    \I__3744\ : InMux
    port map (
            O => \N__16280\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__3743\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16274\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__16274\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0\
        );

    \I__3741\ : InMux
    port map (
            O => \N__16271\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__3740\ : InMux
    port map (
            O => \N__16268\,
            I => \N__16262\
        );

    \I__3739\ : InMux
    port map (
            O => \N__16267\,
            I => \N__16262\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__16262\,
            I => \N__16259\
        );

    \I__3737\ : Span4Mux_v
    port map (
            O => \N__16259\,
            I => \N__16256\
        );

    \I__3736\ : Odrv4
    port map (
            O => \N__16256\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__16253\,
            I => \N__16250\
        );

    \I__3734\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16244\
        );

    \I__3733\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16244\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__16244\,
            I => \N__16240\
        );

    \I__3731\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16237\
        );

    \I__3730\ : Span4Mux_s2_h
    port map (
            O => \N__16240\,
            I => \N__16234\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__16237\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__16234\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__16229\,
            I => \N__16226\
        );

    \I__3726\ : InMux
    port map (
            O => \N__16226\,
            I => \N__16223\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__16223\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6\
        );

    \I__3724\ : InMux
    port map (
            O => \N__16220\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__3723\ : InMux
    port map (
            O => \N__16217\,
            I => \N__16213\
        );

    \I__3722\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16210\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__16213\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__16210\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__16205\,
            I => \N__16202\
        );

    \I__3718\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16199\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__16199\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\
        );

    \I__3716\ : InMux
    port map (
            O => \N__16196\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__3715\ : InMux
    port map (
            O => \N__16193\,
            I => \N__16190\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__16190\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__16187\,
            I => \N__16183\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__16186\,
            I => \N__16180\
        );

    \I__3711\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16175\
        );

    \I__3710\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16175\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__16175\,
            I => charx_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__3708\ : InMux
    port map (
            O => \N__16172\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__3707\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__16166\,
            I => charx_if_generate_plus_mult1_un61_sum_axb_5
        );

    \I__3705\ : InMux
    port map (
            O => \N__16163\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__16160\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_\
        );

    \I__3703\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16152\
        );

    \I__3702\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16149\
        );

    \I__3701\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16146\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__16152\,
            I => \N__16140\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__16149\,
            I => \N__16140\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__16146\,
            I => \N__16137\
        );

    \I__3697\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16132\
        );

    \I__3696\ : Span4Mux_v
    port map (
            O => \N__16140\,
            I => \N__16126\
        );

    \I__3695\ : Span4Mux_v
    port map (
            O => \N__16137\,
            I => \N__16126\
        );

    \I__3694\ : InMux
    port map (
            O => \N__16136\,
            I => \N__16123\
        );

    \I__3693\ : InMux
    port map (
            O => \N__16135\,
            I => \N__16120\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__16132\,
            I => \N__16117\
        );

    \I__3691\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16114\
        );

    \I__3690\ : Sp12to4
    port map (
            O => \N__16126\,
            I => \N__16109\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__16123\,
            I => \N__16109\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__16120\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__16117\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__16114\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__3685\ : Odrv12
    port map (
            O => \N__16109\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__3684\ : InMux
    port map (
            O => \N__16100\,
            I => \N__16097\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__16097\,
            I => charx_if_generate_plus_mult1_un54_sum_i
        );

    \I__3682\ : InMux
    port map (
            O => \N__16094\,
            I => \N__16091\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__16091\,
            I => un5_rowlto2_i
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__16088\,
            I => \N__16075\
        );

    \I__3679\ : CascadeMux
    port map (
            O => \N__16087\,
            I => \N__16072\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__16086\,
            I => \N__16067\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__16085\,
            I => \N__16062\
        );

    \I__3676\ : CascadeMux
    port map (
            O => \N__16084\,
            I => \N__16045\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__16083\,
            I => \N__16042\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__16082\,
            I => \N__16039\
        );

    \I__3673\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16026\
        );

    \I__3672\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16026\
        );

    \I__3671\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16026\
        );

    \I__3670\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16026\
        );

    \I__3669\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16019\
        );

    \I__3668\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16019\
        );

    \I__3667\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16019\
        );

    \I__3666\ : InMux
    port map (
            O => \N__16070\,
            I => \N__16004\
        );

    \I__3665\ : InMux
    port map (
            O => \N__16067\,
            I => \N__16004\
        );

    \I__3664\ : InMux
    port map (
            O => \N__16066\,
            I => \N__15994\
        );

    \I__3663\ : InMux
    port map (
            O => \N__16065\,
            I => \N__15994\
        );

    \I__3662\ : InMux
    port map (
            O => \N__16062\,
            I => \N__15994\
        );

    \I__3661\ : InMux
    port map (
            O => \N__16061\,
            I => \N__15994\
        );

    \I__3660\ : InMux
    port map (
            O => \N__16060\,
            I => \N__15981\
        );

    \I__3659\ : InMux
    port map (
            O => \N__16059\,
            I => \N__15981\
        );

    \I__3658\ : InMux
    port map (
            O => \N__16058\,
            I => \N__15981\
        );

    \I__3657\ : InMux
    port map (
            O => \N__16057\,
            I => \N__15981\
        );

    \I__3656\ : InMux
    port map (
            O => \N__16056\,
            I => \N__15981\
        );

    \I__3655\ : InMux
    port map (
            O => \N__16055\,
            I => \N__15981\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16054\,
            I => \N__15978\
        );

    \I__3653\ : InMux
    port map (
            O => \N__16053\,
            I => \N__15967\
        );

    \I__3652\ : InMux
    port map (
            O => \N__16052\,
            I => \N__15967\
        );

    \I__3651\ : InMux
    port map (
            O => \N__16051\,
            I => \N__15967\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16050\,
            I => \N__15967\
        );

    \I__3649\ : InMux
    port map (
            O => \N__16049\,
            I => \N__15967\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16048\,
            I => \N__15956\
        );

    \I__3647\ : InMux
    port map (
            O => \N__16045\,
            I => \N__15956\
        );

    \I__3646\ : InMux
    port map (
            O => \N__16042\,
            I => \N__15956\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16039\,
            I => \N__15956\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16038\,
            I => \N__15956\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16037\,
            I => \N__15949\
        );

    \I__3642\ : InMux
    port map (
            O => \N__16036\,
            I => \N__15949\
        );

    \I__3641\ : InMux
    port map (
            O => \N__16035\,
            I => \N__15949\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__16026\,
            I => \N__15946\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16019\,
            I => \N__15943\
        );

    \I__3638\ : InMux
    port map (
            O => \N__16018\,
            I => \N__15936\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16017\,
            I => \N__15936\
        );

    \I__3636\ : InMux
    port map (
            O => \N__16016\,
            I => \N__15936\
        );

    \I__3635\ : InMux
    port map (
            O => \N__16015\,
            I => \N__15933\
        );

    \I__3634\ : InMux
    port map (
            O => \N__16014\,
            I => \N__15930\
        );

    \I__3633\ : InMux
    port map (
            O => \N__16013\,
            I => \N__15923\
        );

    \I__3632\ : InMux
    port map (
            O => \N__16012\,
            I => \N__15923\
        );

    \I__3631\ : InMux
    port map (
            O => \N__16011\,
            I => \N__15923\
        );

    \I__3630\ : InMux
    port map (
            O => \N__16010\,
            I => \N__15918\
        );

    \I__3629\ : InMux
    port map (
            O => \N__16009\,
            I => \N__15918\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__16004\,
            I => \N__15915\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16003\,
            I => \N__15912\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__15994\,
            I => \N__15907\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__15981\,
            I => \N__15907\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__15978\,
            I => \N__15894\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__15967\,
            I => \N__15894\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__15956\,
            I => \N__15894\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15894\
        );

    \I__3620\ : Span4Mux_s3_v
    port map (
            O => \N__15946\,
            I => \N__15894\
        );

    \I__3619\ : Span4Mux_s3_v
    port map (
            O => \N__15943\,
            I => \N__15894\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__15936\,
            I => un5_rowlto2
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__15933\,
            I => un5_rowlto2
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__15930\,
            I => un5_rowlto2
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__15923\,
            I => un5_rowlto2
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__15918\,
            I => un5_rowlto2
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__15915\,
            I => un5_rowlto2
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__15912\,
            I => un5_rowlto2
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__15907\,
            I => un5_rowlto2
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__15894\,
            I => un5_rowlto2
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__15875\,
            I => \N__15870\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__15874\,
            I => \N__15865\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__15873\,
            I => \N__15859\
        );

    \I__3606\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15843\
        );

    \I__3605\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15843\
        );

    \I__3604\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15836\
        );

    \I__3603\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15836\
        );

    \I__3602\ : CascadeMux
    port map (
            O => \N__15864\,
            I => \N__15832\
        );

    \I__3601\ : CascadeMux
    port map (
            O => \N__15863\,
            I => \N__15829\
        );

    \I__3600\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15825\
        );

    \I__3599\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15822\
        );

    \I__3598\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15817\
        );

    \I__3597\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15817\
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__15856\,
            I => \N__15814\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \N__15808\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__15854\,
            I => \N__15803\
        );

    \I__3593\ : CascadeMux
    port map (
            O => \N__15853\,
            I => \N__15800\
        );

    \I__3592\ : CascadeMux
    port map (
            O => \N__15852\,
            I => \N__15795\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__15851\,
            I => \N__15790\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__15850\,
            I => \N__15784\
        );

    \I__3589\ : CascadeMux
    port map (
            O => \N__15849\,
            I => \N__15781\
        );

    \I__3588\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15778\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__15843\,
            I => \N__15775\
        );

    \I__3586\ : InMux
    port map (
            O => \N__15842\,
            I => \N__15770\
        );

    \I__3585\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15770\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__15836\,
            I => \N__15767\
        );

    \I__3583\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15758\
        );

    \I__3582\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15758\
        );

    \I__3581\ : InMux
    port map (
            O => \N__15829\,
            I => \N__15758\
        );

    \I__3580\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15758\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__15825\,
            I => \N__15751\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__15822\,
            I => \N__15751\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__15817\,
            I => \N__15751\
        );

    \I__3576\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15740\
        );

    \I__3575\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15740\
        );

    \I__3574\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15740\
        );

    \I__3573\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15740\
        );

    \I__3572\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15740\
        );

    \I__3571\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15729\
        );

    \I__3570\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15729\
        );

    \I__3569\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15729\
        );

    \I__3568\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15729\
        );

    \I__3567\ : InMux
    port map (
            O => \N__15799\,
            I => \N__15729\
        );

    \I__3566\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15718\
        );

    \I__3565\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15718\
        );

    \I__3564\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15718\
        );

    \I__3563\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15718\
        );

    \I__3562\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15718\
        );

    \I__3561\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15707\
        );

    \I__3560\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15707\
        );

    \I__3559\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15707\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15707\
        );

    \I__3557\ : InMux
    port map (
            O => \N__15781\,
            I => \N__15707\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__15778\,
            I => un5_rowlto0
        );

    \I__3555\ : Odrv12
    port map (
            O => \N__15775\,
            I => un5_rowlto0
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__15770\,
            I => un5_rowlto0
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__15767\,
            I => un5_rowlto0
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__15758\,
            I => un5_rowlto0
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__15751\,
            I => un5_rowlto0
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__15740\,
            I => un5_rowlto0
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__15729\,
            I => un5_rowlto0
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__15718\,
            I => un5_rowlto0
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__15707\,
            I => un5_rowlto0
        );

    \I__3546\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15670\
        );

    \I__3545\ : InMux
    port map (
            O => \N__15685\,
            I => \N__15667\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__15684\,
            I => \N__15650\
        );

    \I__3543\ : InMux
    port map (
            O => \N__15683\,
            I => \N__15645\
        );

    \I__3542\ : InMux
    port map (
            O => \N__15682\,
            I => \N__15645\
        );

    \I__3541\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15640\
        );

    \I__3540\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15640\
        );

    \I__3539\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15633\
        );

    \I__3538\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15633\
        );

    \I__3537\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15633\
        );

    \I__3536\ : CascadeMux
    port map (
            O => \N__15676\,
            I => \N__15628\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__15675\,
            I => \N__15625\
        );

    \I__3534\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15619\
        );

    \I__3533\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15619\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__15670\,
            I => \N__15614\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__15667\,
            I => \N__15614\
        );

    \I__3530\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15609\
        );

    \I__3529\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15609\
        );

    \I__3528\ : InMux
    port map (
            O => \N__15664\,
            I => \N__15598\
        );

    \I__3527\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15598\
        );

    \I__3526\ : InMux
    port map (
            O => \N__15662\,
            I => \N__15598\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15661\,
            I => \N__15598\
        );

    \I__3524\ : InMux
    port map (
            O => \N__15660\,
            I => \N__15598\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__15659\,
            I => \N__15595\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__15658\,
            I => \N__15590\
        );

    \I__3521\ : CascadeMux
    port map (
            O => \N__15657\,
            I => \N__15584\
        );

    \I__3520\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15571\
        );

    \I__3519\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15571\
        );

    \I__3518\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15571\
        );

    \I__3517\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15571\
        );

    \I__3516\ : InMux
    port map (
            O => \N__15650\,
            I => \N__15571\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__15645\,
            I => \N__15568\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__15640\,
            I => \N__15563\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__15633\,
            I => \N__15563\
        );

    \I__3512\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15560\
        );

    \I__3511\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15551\
        );

    \I__3510\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15551\
        );

    \I__3509\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15551\
        );

    \I__3508\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15551\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__15619\,
            I => \N__15542\
        );

    \I__3506\ : Span4Mux_v
    port map (
            O => \N__15614\,
            I => \N__15542\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__15609\,
            I => \N__15542\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__15598\,
            I => \N__15542\
        );

    \I__3503\ : InMux
    port map (
            O => \N__15595\,
            I => \N__15533\
        );

    \I__3502\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15533\
        );

    \I__3501\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15533\
        );

    \I__3500\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15533\
        );

    \I__3499\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15526\
        );

    \I__3498\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15526\
        );

    \I__3497\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15526\
        );

    \I__3496\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15519\
        );

    \I__3495\ : InMux
    port map (
            O => \N__15583\,
            I => \N__15519\
        );

    \I__3494\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15519\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__15571\,
            I => un5_rowlto1
        );

    \I__3492\ : Odrv12
    port map (
            O => \N__15568\,
            I => un5_rowlto1
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__15563\,
            I => un5_rowlto1
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15560\,
            I => un5_rowlto1
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__15551\,
            I => un5_rowlto1
        );

    \I__3488\ : Odrv4
    port map (
            O => \N__15542\,
            I => un5_rowlto1
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__15533\,
            I => un5_rowlto1
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__15526\,
            I => un5_rowlto1
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__15519\,
            I => un5_rowlto1
        );

    \I__3484\ : InMux
    port map (
            O => \N__15500\,
            I => \N__15482\
        );

    \I__3483\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15482\
        );

    \I__3482\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15482\
        );

    \I__3481\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15482\
        );

    \I__3480\ : InMux
    port map (
            O => \N__15496\,
            I => \N__15462\
        );

    \I__3479\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15462\
        );

    \I__3478\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15453\
        );

    \I__3477\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15453\
        );

    \I__3476\ : InMux
    port map (
            O => \N__15492\,
            I => \N__15453\
        );

    \I__3475\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15453\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__15482\,
            I => \N__15450\
        );

    \I__3473\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15439\
        );

    \I__3472\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15439\
        );

    \I__3471\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15439\
        );

    \I__3470\ : InMux
    port map (
            O => \N__15478\,
            I => \N__15439\
        );

    \I__3469\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15439\
        );

    \I__3468\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15434\
        );

    \I__3467\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15434\
        );

    \I__3466\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15427\
        );

    \I__3465\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15427\
        );

    \I__3464\ : InMux
    port map (
            O => \N__15472\,
            I => \N__15427\
        );

    \I__3463\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15420\
        );

    \I__3462\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15420\
        );

    \I__3461\ : InMux
    port map (
            O => \N__15469\,
            I => \N__15420\
        );

    \I__3460\ : InMux
    port map (
            O => \N__15468\,
            I => \N__15415\
        );

    \I__3459\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15415\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__15462\,
            I => \N__15406\
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__15453\,
            I => \N__15406\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__15450\,
            I => \N__15403\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__15439\,
            I => \N__15396\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__15434\,
            I => \N__15396\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__15427\,
            I => \N__15396\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__15420\,
            I => \N__15391\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__15415\,
            I => \N__15391\
        );

    \I__3450\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15386\
        );

    \I__3449\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15386\
        );

    \I__3448\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15378\
        );

    \I__3447\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15378\
        );

    \I__3446\ : Span4Mux_v
    port map (
            O => \N__15406\,
            I => \N__15373\
        );

    \I__3445\ : Span4Mux_v
    port map (
            O => \N__15403\,
            I => \N__15373\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__15396\,
            I => \N__15366\
        );

    \I__3443\ : Span4Mux_v
    port map (
            O => \N__15391\,
            I => \N__15366\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__15386\,
            I => \N__15366\
        );

    \I__3441\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15363\
        );

    \I__3440\ : InMux
    port map (
            O => \N__15384\,
            I => \N__15358\
        );

    \I__3439\ : InMux
    port map (
            O => \N__15383\,
            I => \N__15358\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__15378\,
            I => un5_rowlto3
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__15373\,
            I => un5_rowlto3
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__15366\,
            I => un5_rowlto3
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__15363\,
            I => un5_rowlto3
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__15358\,
            I => un5_rowlto3
        );

    \I__3433\ : InMux
    port map (
            O => \N__15347\,
            I => \N__15344\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__15344\,
            I => \un116_pixel_2_amZ0Z_1\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \N__15338\
        );

    \I__3430\ : InMux
    port map (
            O => \N__15338\,
            I => \N__15335\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__15335\,
            I => \N__15332\
        );

    \I__3428\ : Span4Mux_s2_h
    port map (
            O => \N__15332\,
            I => \N__15329\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__15329\,
            I => charx_if_generate_plus_mult1_un47_sum_i_5
        );

    \I__3426\ : InMux
    port map (
            O => \N__15326\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__3425\ : InMux
    port map (
            O => \N__15323\,
            I => \N__15320\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__3423\ : Span4Mux_s2_h
    port map (
            O => \N__15317\,
            I => \N__15314\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__15314\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\
        );

    \I__3421\ : InMux
    port map (
            O => \N__15311\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__3420\ : InMux
    port map (
            O => \N__15308\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__3419\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15302\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__15302\,
            I => \N__15299\
        );

    \I__3417\ : Span4Mux_v
    port map (
            O => \N__15299\,
            I => \N__15296\
        );

    \I__3416\ : Odrv4
    port map (
            O => \N__15296\,
            I => charx_if_generate_plus_mult1_un54_sum_axb_5
        );

    \I__3415\ : InMux
    port map (
            O => \N__15293\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__15290\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7_cascade_\
        );

    \I__3413\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15281\
        );

    \I__3412\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15276\
        );

    \I__3411\ : InMux
    port map (
            O => \N__15285\,
            I => \N__15273\
        );

    \I__3410\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15270\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__15281\,
            I => \N__15267\
        );

    \I__3408\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15264\
        );

    \I__3407\ : InMux
    port map (
            O => \N__15279\,
            I => \N__15261\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__15276\,
            I => \N__15256\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__15273\,
            I => \N__15256\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__15270\,
            I => \N__15253\
        );

    \I__3403\ : Span4Mux_h
    port map (
            O => \N__15267\,
            I => \N__15250\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__15264\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__15261\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__15256\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__3399\ : Odrv12
    port map (
            O => \N__15253\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__15250\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__3397\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__15236\,
            I => charx_if_generate_plus_mult1_un47_sum_i
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__3394\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__15227\,
            I => \N__15224\
        );

    \I__3392\ : Span4Mux_h
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__15221\,
            I => \N_302_i_0\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__15218\,
            I => \beamY_RNITQPUS72Z0Z_0_cascade_\
        );

    \I__3389\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15212\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__15212\,
            I => un116_pixel_3_1_0
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \N__15206\
        );

    \I__3386\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__15203\,
            I => \beamY_RNI6B7UAL1Z0Z_1\
        );

    \I__3384\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15197\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__15197\,
            I => \N__15194\
        );

    \I__3382\ : Span4Mux_h
    port map (
            O => \N__15194\,
            I => \N__15190\
        );

    \I__3381\ : InMux
    port map (
            O => \N__15193\,
            I => \N__15187\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__15190\,
            I => m31
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__15187\,
            I => m31
        );

    \I__3378\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15179\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__15179\,
            I => \un116_pixel_4_1Z0Z_0\
        );

    \I__3376\ : InMux
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__15173\,
            I => m38
        );

    \I__3374\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15167\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15157\
        );

    \I__3372\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15154\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__15165\,
            I => \N__15150\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__15164\,
            I => \N__15147\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__15163\,
            I => \N__15139\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__15162\,
            I => \N__15134\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__15161\,
            I => \N__15129\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__15160\,
            I => \N__15124\
        );

    \I__3365\ : Span4Mux_h
    port map (
            O => \N__15157\,
            I => \N__15119\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__15154\,
            I => \N__15119\
        );

    \I__3363\ : InMux
    port map (
            O => \N__15153\,
            I => \N__15110\
        );

    \I__3362\ : InMux
    port map (
            O => \N__15150\,
            I => \N__15110\
        );

    \I__3361\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15110\
        );

    \I__3360\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15110\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__15145\,
            I => \N__15103\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__15144\,
            I => \N__15098\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__15143\,
            I => \N__15094\
        );

    \I__3356\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15091\
        );

    \I__3355\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15088\
        );

    \I__3354\ : InMux
    port map (
            O => \N__15138\,
            I => \N__15085\
        );

    \I__3353\ : InMux
    port map (
            O => \N__15137\,
            I => \N__15082\
        );

    \I__3352\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15079\
        );

    \I__3351\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15076\
        );

    \I__3350\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15073\
        );

    \I__3349\ : InMux
    port map (
            O => \N__15129\,
            I => \N__15066\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15066\
        );

    \I__3347\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15066\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15063\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__15119\,
            I => \N__15058\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__15110\,
            I => \N__15058\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15109\,
            I => \N__15053\
        );

    \I__3342\ : InMux
    port map (
            O => \N__15108\,
            I => \N__15053\
        );

    \I__3341\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15049\
        );

    \I__3340\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15038\
        );

    \I__3339\ : InMux
    port map (
            O => \N__15103\,
            I => \N__15038\
        );

    \I__3338\ : InMux
    port map (
            O => \N__15102\,
            I => \N__15038\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15101\,
            I => \N__15038\
        );

    \I__3336\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15038\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__15097\,
            I => \N__15032\
        );

    \I__3334\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15029\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__15091\,
            I => \N__15026\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__15088\,
            I => \N__15019\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__15085\,
            I => \N__15019\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__15082\,
            I => \N__15019\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__15079\,
            I => \N__15016\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__15076\,
            I => \N__15013\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__15073\,
            I => \N__15010\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__15066\,
            I => \N__15001\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__15063\,
            I => \N__15001\
        );

    \I__3324\ : Span4Mux_v
    port map (
            O => \N__15058\,
            I => \N__15001\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__15053\,
            I => \N__15001\
        );

    \I__3322\ : InMux
    port map (
            O => \N__15052\,
            I => \N__14997\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__15049\,
            I => \N__14994\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__15038\,
            I => \N__14991\
        );

    \I__3319\ : InMux
    port map (
            O => \N__15037\,
            I => \N__14988\
        );

    \I__3318\ : InMux
    port map (
            O => \N__15036\,
            I => \N__14981\
        );

    \I__3317\ : InMux
    port map (
            O => \N__15035\,
            I => \N__14981\
        );

    \I__3316\ : InMux
    port map (
            O => \N__15032\,
            I => \N__14981\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__15029\,
            I => \N__14974\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__15026\,
            I => \N__14974\
        );

    \I__3313\ : Span4Mux_h
    port map (
            O => \N__15019\,
            I => \N__14974\
        );

    \I__3312\ : Span4Mux_h
    port map (
            O => \N__15016\,
            I => \N__14969\
        );

    \I__3311\ : Span4Mux_h
    port map (
            O => \N__15013\,
            I => \N__14969\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__15010\,
            I => \N__14964\
        );

    \I__3309\ : Span4Mux_h
    port map (
            O => \N__15001\,
            I => \N__14964\
        );

    \I__3308\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14961\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__14997\,
            I => \beamYZ0Z_0\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__14994\,
            I => \beamYZ0Z_0\
        );

    \I__3305\ : Odrv4
    port map (
            O => \N__14991\,
            I => \beamYZ0Z_0\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__14988\,
            I => \beamYZ0Z_0\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__14981\,
            I => \beamYZ0Z_0\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__14974\,
            I => \beamYZ0Z_0\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__14969\,
            I => \beamYZ0Z_0\
        );

    \I__3300\ : Odrv4
    port map (
            O => \N__14964\,
            I => \beamYZ0Z_0\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__14961\,
            I => \beamYZ0Z_0\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__14942\,
            I => \m38_cascade_\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__14939\,
            I => \N__14931\
        );

    \I__3296\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14926\
        );

    \I__3295\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14917\
        );

    \I__3294\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14914\
        );

    \I__3293\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14909\
        );

    \I__3292\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14909\
        );

    \I__3291\ : InMux
    port map (
            O => \N__14931\,
            I => \N__14902\
        );

    \I__3290\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14899\
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__14929\,
            I => \N__14895\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__14926\,
            I => \N__14892\
        );

    \I__3287\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14889\
        );

    \I__3286\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14886\
        );

    \I__3285\ : InMux
    port map (
            O => \N__14923\,
            I => \N__14883\
        );

    \I__3284\ : InMux
    port map (
            O => \N__14922\,
            I => \N__14880\
        );

    \I__3283\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14877\
        );

    \I__3282\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14874\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__14917\,
            I => \N__14870\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__14914\,
            I => \N__14865\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__14909\,
            I => \N__14865\
        );

    \I__3278\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14862\
        );

    \I__3277\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14859\
        );

    \I__3276\ : InMux
    port map (
            O => \N__14906\,
            I => \N__14856\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__14905\,
            I => \N__14851\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__14902\,
            I => \N__14844\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__14899\,
            I => \N__14841\
        );

    \I__3272\ : CascadeMux
    port map (
            O => \N__14898\,
            I => \N__14838\
        );

    \I__3271\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14835\
        );

    \I__3270\ : Span4Mux_v
    port map (
            O => \N__14892\,
            I => \N__14832\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__14889\,
            I => \N__14825\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__14886\,
            I => \N__14825\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__14883\,
            I => \N__14825\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__14880\,
            I => \N__14820\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__14877\,
            I => \N__14820\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__14874\,
            I => \N__14817\
        );

    \I__3263\ : InMux
    port map (
            O => \N__14873\,
            I => \N__14814\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__14870\,
            I => \N__14803\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__14865\,
            I => \N__14803\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__14862\,
            I => \N__14803\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__14859\,
            I => \N__14803\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__14856\,
            I => \N__14803\
        );

    \I__3257\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14800\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14854\,
            I => \N__14797\
        );

    \I__3255\ : InMux
    port map (
            O => \N__14851\,
            I => \N__14794\
        );

    \I__3254\ : InMux
    port map (
            O => \N__14850\,
            I => \N__14787\
        );

    \I__3253\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14787\
        );

    \I__3252\ : InMux
    port map (
            O => \N__14848\,
            I => \N__14787\
        );

    \I__3251\ : InMux
    port map (
            O => \N__14847\,
            I => \N__14784\
        );

    \I__3250\ : Span4Mux_h
    port map (
            O => \N__14844\,
            I => \N__14779\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__14841\,
            I => \N__14779\
        );

    \I__3248\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14776\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__14835\,
            I => \N__14769\
        );

    \I__3246\ : Span4Mux_s2_h
    port map (
            O => \N__14832\,
            I => \N__14769\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__14825\,
            I => \N__14769\
        );

    \I__3244\ : Span4Mux_h
    port map (
            O => \N__14820\,
            I => \N__14760\
        );

    \I__3243\ : Span4Mux_h
    port map (
            O => \N__14817\,
            I => \N__14760\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__14814\,
            I => \N__14760\
        );

    \I__3241\ : Span4Mux_v
    port map (
            O => \N__14803\,
            I => \N__14760\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__14800\,
            I => \beamYZ0Z_1\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__14797\,
            I => \beamYZ0Z_1\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__14794\,
            I => \beamYZ0Z_1\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__14787\,
            I => \beamYZ0Z_1\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__14784\,
            I => \beamYZ0Z_1\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__14779\,
            I => \beamYZ0Z_1\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__14776\,
            I => \beamYZ0Z_1\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__14769\,
            I => \beamYZ0Z_1\
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__14760\,
            I => \beamYZ0Z_1\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__14741\,
            I => \un116_pixel_6_1_1_cascade_\
        );

    \I__3230\ : InMux
    port map (
            O => \N__14738\,
            I => \N__14735\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__14732\,
            I => \N_17\
        );

    \I__3227\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14719\
        );

    \I__3225\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14714\
        );

    \I__3224\ : InMux
    port map (
            O => \N__14724\,
            I => \N__14714\
        );

    \I__3223\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14711\
        );

    \I__3222\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14708\
        );

    \I__3221\ : Span4Mux_h
    port map (
            O => \N__14719\,
            I => \N__14703\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__14714\,
            I => \N__14703\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__14711\,
            I => \N__14700\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__14708\,
            I => \N_321\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__14703\,
            I => \N_321\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__14700\,
            I => \N_321\
        );

    \I__3215\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__14690\,
            I => \un116_pixel_2_bmZ0Z_1\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__14687\,
            I => \beamY_RNI4NRC8D1Z0Z_0_cascade_\
        );

    \I__3212\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14681\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__14681\,
            I => \beamY_RNII25UDD3Z0Z_0\
        );

    \I__3210\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14675\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__14675\,
            I => \N_14\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__14672\,
            I => \un116_pixel_2_ns_1_6_cascade_\
        );

    \I__3207\ : InMux
    port map (
            O => \N__14669\,
            I => \N__14666\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__14666\,
            I => \beamY_RNIH01F2SZ0Z_0\
        );

    \I__3205\ : InMux
    port map (
            O => \N__14663\,
            I => \N__14660\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__14660\,
            I => \un116_pixel_2_ns_1Z0Z_5\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \N_276_0_cascade_\
        );

    \I__3202\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14651\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__14651\,
            I => \N__14648\
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__14648\,
            I => \beamY_RNII25UDD3_3Z0Z_0\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14642\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__14642\,
            I => m7
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__14639\,
            I => \m7_cascade_\
        );

    \I__3196\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14633\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__14633\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3\
        );

    \I__3194\ : InMux
    port map (
            O => \N__14630\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__3192\ : InMux
    port map (
            O => \N__14624\,
            I => \N__14621\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__14621\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0\
        );

    \I__3190\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14609\
        );

    \I__3189\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14609\
        );

    \I__3188\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14609\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__14609\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\
        );

    \I__3186\ : InMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__14603\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__14600\,
            I => \N__14596\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__14599\,
            I => \N__14593\
        );

    \I__3182\ : InMux
    port map (
            O => \N__14596\,
            I => \N__14588\
        );

    \I__3181\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14588\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__14588\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\
        );

    \I__3179\ : InMux
    port map (
            O => \N__14585\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4
        );

    \I__3178\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14575\
        );

    \I__3177\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14572\
        );

    \I__3176\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14565\
        );

    \I__3175\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14565\
        );

    \I__3174\ : InMux
    port map (
            O => \N__14578\,
            I => \N__14565\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__14575\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__14572\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__14565\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\
        );

    \I__3170\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14555\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__14555\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPBZ0Z3\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__14552\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_\
        );

    \I__3167\ : CascadeMux
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__3166\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14540\
        );

    \I__3165\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14540\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__14540\,
            I => \un114_pixel_6_1_5__font_un126_pixel_m_1Z0Z_1\
        );

    \I__3163\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14528\
        );

    \I__3162\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14525\
        );

    \I__3161\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14518\
        );

    \I__3160\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14518\
        );

    \I__3159\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14518\
        );

    \I__3158\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14513\
        );

    \I__3157\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14513\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__14528\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__14525\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__14518\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__14513\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__3152\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14494\
        );

    \I__3151\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14487\
        );

    \I__3150\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14487\
        );

    \I__3149\ : InMux
    port map (
            O => \N__14501\,
            I => \N__14487\
        );

    \I__3148\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14484\
        );

    \I__3147\ : InMux
    port map (
            O => \N__14499\,
            I => \N__14481\
        );

    \I__3146\ : InMux
    port map (
            O => \N__14498\,
            I => \N__14478\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__14497\,
            I => \N__14471\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__14494\,
            I => \N__14466\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__14487\,
            I => \N__14466\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__14484\,
            I => \N__14461\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__14481\,
            I => \N__14461\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__14478\,
            I => \N__14458\
        );

    \I__3139\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14455\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__14476\,
            I => \N__14452\
        );

    \I__3137\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14447\
        );

    \I__3136\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14447\
        );

    \I__3135\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14444\
        );

    \I__3134\ : Span12Mux_s6_h
    port map (
            O => \N__14466\,
            I => \N__14441\
        );

    \I__3133\ : Span4Mux_v
    port map (
            O => \N__14461\,
            I => \N__14438\
        );

    \I__3132\ : Span12Mux_s10_v
    port map (
            O => \N__14458\,
            I => \N__14435\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__14455\,
            I => \N__14432\
        );

    \I__3130\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14429\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__14447\,
            I => \beamXZ0Z_0\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__14444\,
            I => \beamXZ0Z_0\
        );

    \I__3127\ : Odrv12
    port map (
            O => \N__14441\,
            I => \beamXZ0Z_0\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__14438\,
            I => \beamXZ0Z_0\
        );

    \I__3125\ : Odrv12
    port map (
            O => \N__14435\,
            I => \beamXZ0Z_0\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__14432\,
            I => \beamXZ0Z_0\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__14429\,
            I => \beamXZ0Z_0\
        );

    \I__3122\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14409\
        );

    \I__3121\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14406\
        );

    \I__3120\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14403\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__14409\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__14406\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__14403\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__14396\,
            I => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\
        );

    \I__3115\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14390\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__14390\,
            I => \un114_pixel_6_1_5__font_un126_pixel_m_1_1Z0Z_1\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__14387\,
            I => \m15_cascade_\
        );

    \I__3112\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14377\
        );

    \I__3111\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14372\
        );

    \I__3110\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14372\
        );

    \I__3109\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14369\
        );

    \I__3108\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14366\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__14377\,
            I => \N__14363\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__14372\,
            I => \N__14360\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__14369\,
            I => \un114_pixel_0_1__N_6_mux\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__14366\,
            I => \un114_pixel_0_1__N_6_mux\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__14363\,
            I => \un114_pixel_0_1__N_6_mux\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__14360\,
            I => \un114_pixel_0_1__N_6_mux\
        );

    \I__3101\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14347\
        );

    \I__3100\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14342\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__14347\,
            I => \N__14339\
        );

    \I__3098\ : InMux
    port map (
            O => \N__14346\,
            I => \N__14336\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__14345\,
            I => \N__14331\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14326\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__14339\,
            I => \N__14321\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__14336\,
            I => \N__14321\
        );

    \I__3093\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14316\
        );

    \I__3092\ : InMux
    port map (
            O => \N__14334\,
            I => \N__14316\
        );

    \I__3091\ : InMux
    port map (
            O => \N__14331\,
            I => \N__14313\
        );

    \I__3090\ : InMux
    port map (
            O => \N__14330\,
            I => \N__14310\
        );

    \I__3089\ : InMux
    port map (
            O => \N__14329\,
            I => \N__14307\
        );

    \I__3088\ : Span4Mux_h
    port map (
            O => \N__14326\,
            I => \N__14304\
        );

    \I__3087\ : Span4Mux_h
    port map (
            O => \N__14321\,
            I => \N__14301\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__14316\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__14313\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__14310\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__14307\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__14304\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__14301\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__3080\ : InMux
    port map (
            O => \N__14288\,
            I => \N__14285\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__14285\,
            I => charx_if_generate_plus_mult1_un40_sum_i
        );

    \I__3078\ : InMux
    port map (
            O => \N__14282\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1
        );

    \I__3077\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14267\
        );

    \I__3076\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14262\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__14277\,
            I => \N__14259\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__14276\,
            I => \N__14256\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__14275\,
            I => \N__14253\
        );

    \I__3072\ : InMux
    port map (
            O => \N__14274\,
            I => \N__14247\
        );

    \I__3071\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14242\
        );

    \I__3070\ : InMux
    port map (
            O => \N__14272\,
            I => \N__14242\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__14271\,
            I => \N__14239\
        );

    \I__3068\ : InMux
    port map (
            O => \N__14270\,
            I => \N__14233\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__14267\,
            I => \N__14230\
        );

    \I__3066\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14227\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__14265\,
            I => \N__14223\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__14262\,
            I => \N__14218\
        );

    \I__3063\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14215\
        );

    \I__3062\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14210\
        );

    \I__3061\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14210\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__14252\,
            I => \N__14207\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__14251\,
            I => \N__14204\
        );

    \I__3058\ : IoInMux
    port map (
            O => \N__14250\,
            I => \N__14201\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__14247\,
            I => \N__14196\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__14242\,
            I => \N__14196\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14191\
        );

    \I__3054\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14191\
        );

    \I__3053\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14188\
        );

    \I__3052\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14185\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__14233\,
            I => \N__14181\
        );

    \I__3050\ : Span4Mux_v
    port map (
            O => \N__14230\,
            I => \N__14176\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__14227\,
            I => \N__14176\
        );

    \I__3048\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14173\
        );

    \I__3047\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14168\
        );

    \I__3046\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14168\
        );

    \I__3045\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14165\
        );

    \I__3044\ : Span4Mux_v
    port map (
            O => \N__14218\,
            I => \N__14158\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__14215\,
            I => \N__14158\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__14210\,
            I => \N__14158\
        );

    \I__3041\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14155\
        );

    \I__3040\ : InMux
    port map (
            O => \N__14204\,
            I => \N__14152\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__14201\,
            I => \N__14149\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__14196\,
            I => \N__14140\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__14191\,
            I => \N__14140\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__14188\,
            I => \N__14140\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__14185\,
            I => \N__14140\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14137\
        );

    \I__3033\ : Span4Mux_v
    port map (
            O => \N__14181\,
            I => \N__14126\
        );

    \I__3032\ : Span4Mux_h
    port map (
            O => \N__14176\,
            I => \N__14126\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__14173\,
            I => \N__14126\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__14168\,
            I => \N__14126\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__14165\,
            I => \N__14126\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__14158\,
            I => \N__14119\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__14155\,
            I => \N__14119\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__14152\,
            I => \N__14119\
        );

    \I__3025\ : IoSpan4Mux
    port map (
            O => \N__14149\,
            I => \N__14116\
        );

    \I__3024\ : Span4Mux_h
    port map (
            O => \N__14140\,
            I => \N__14111\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__14137\,
            I => \N__14111\
        );

    \I__3022\ : Span4Mux_v
    port map (
            O => \N__14126\,
            I => \N__14108\
        );

    \I__3021\ : Span4Mux_h
    port map (
            O => \N__14119\,
            I => \N__14103\
        );

    \I__3020\ : Span4Mux_s1_v
    port map (
            O => \N__14116\,
            I => \N__14103\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__14111\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__14108\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__14103\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3016\ : InMux
    port map (
            O => \N__14096\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2
        );

    \I__3015\ : InMux
    port map (
            O => \N__14093\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3
        );

    \I__3014\ : InMux
    port map (
            O => \N__14090\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4
        );

    \I__3013\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14084\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__14084\,
            I => \N__14081\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__14081\,
            I => \un114_pixel_6_1_5__g2_0_1\
        );

    \I__3010\ : InMux
    port map (
            O => \N__14078\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1
        );

    \I__3009\ : CascadeMux
    port map (
            O => \N__14075\,
            I => \N__14071\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__14074\,
            I => \N__14068\
        );

    \I__3007\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14063\
        );

    \I__3006\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14063\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__14063\,
            I => charx_if_generate_plus_mult1_un33_sum_i_5
        );

    \I__3004\ : InMux
    port map (
            O => \N__14060\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__3003\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14054\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__14054\,
            I => charx_if_generate_plus_mult1_un40_sum_axb_5
        );

    \I__3001\ : InMux
    port map (
            O => \N__14051\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__3000\ : InMux
    port map (
            O => \N__14048\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_1
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__14045\,
            I => \N__14042\
        );

    \I__2998\ : InMux
    port map (
            O => \N__14042\,
            I => \N__14039\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__14039\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\
        );

    \I__2996\ : InMux
    port map (
            O => \N__14036\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__2995\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14030\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__14030\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\
        );

    \I__2993\ : InMux
    port map (
            O => \N__14027\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__2992\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14021\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__14021\,
            I => charx_if_generate_plus_mult1_un47_sum_axb_5
        );

    \I__2990\ : InMux
    port map (
            O => \N__14018\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__14015\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_\
        );

    \I__2988\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14007\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14011\,
            I => \N__14002\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14010\,
            I => \N__14002\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__14007\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__14002\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__13997\,
            I => \N__13993\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__2981\ : InMux
    port map (
            O => \N__13993\,
            I => \N__13985\
        );

    \I__2980\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13985\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__13985\,
            I => charx_if_generate_plus_mult1_un40_sum_i_5
        );

    \I__2978\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__13979\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\
        );

    \I__2976\ : InMux
    port map (
            O => \N__13976\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__2974\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__13967\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\
        );

    \I__2972\ : InMux
    port map (
            O => \N__13964\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__13961\,
            I => \N__13949\
        );

    \I__2970\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13940\
        );

    \I__2969\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13940\
        );

    \I__2968\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13937\
        );

    \I__2967\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13934\
        );

    \I__2966\ : InMux
    port map (
            O => \N__13956\,
            I => \N__13931\
        );

    \I__2965\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13922\
        );

    \I__2964\ : InMux
    port map (
            O => \N__13954\,
            I => \N__13922\
        );

    \I__2963\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13922\
        );

    \I__2962\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13922\
        );

    \I__2961\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13919\
        );

    \I__2960\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13909\
        );

    \I__2959\ : InMux
    port map (
            O => \N__13947\,
            I => \N__13909\
        );

    \I__2958\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13909\
        );

    \I__2957\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13909\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__13940\,
            I => \N__13906\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__13937\,
            I => \N__13901\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__13934\,
            I => \N__13901\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__13931\,
            I => \N__13894\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__13922\,
            I => \N__13894\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__13919\,
            I => \N__13894\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__13918\,
            I => \N__13883\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__13909\,
            I => \N__13880\
        );

    \I__2948\ : Span4Mux_v
    port map (
            O => \N__13906\,
            I => \N__13875\
        );

    \I__2947\ : Span4Mux_v
    port map (
            O => \N__13901\,
            I => \N__13875\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__13894\,
            I => \N__13872\
        );

    \I__2945\ : InMux
    port map (
            O => \N__13893\,
            I => \N__13857\
        );

    \I__2944\ : InMux
    port map (
            O => \N__13892\,
            I => \N__13857\
        );

    \I__2943\ : InMux
    port map (
            O => \N__13891\,
            I => \N__13857\
        );

    \I__2942\ : InMux
    port map (
            O => \N__13890\,
            I => \N__13857\
        );

    \I__2941\ : InMux
    port map (
            O => \N__13889\,
            I => \N__13857\
        );

    \I__2940\ : InMux
    port map (
            O => \N__13888\,
            I => \N__13857\
        );

    \I__2939\ : InMux
    port map (
            O => \N__13887\,
            I => \N__13857\
        );

    \I__2938\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13852\
        );

    \I__2937\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13852\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__13880\,
            I => \CO3_0\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__13875\,
            I => \CO3_0\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__13872\,
            I => \CO3_0\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__13857\,
            I => \CO3_0\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__13852\,
            I => \CO3_0\
        );

    \I__2931\ : InMux
    port map (
            O => \N__13841\,
            I => \N__13838\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__13838\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\
        );

    \I__2929\ : InMux
    port map (
            O => \N__13835\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__13832\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0_cascade_\
        );

    \I__2927\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13820\
        );

    \I__2926\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13820\
        );

    \I__2925\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13820\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__13820\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__13817\,
            I => \N__13813\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__13816\,
            I => \N__13810\
        );

    \I__2921\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13805\
        );

    \I__2920\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13805\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__13805\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\
        );

    \I__2918\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13799\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__13799\,
            I => \N__13796\
        );

    \I__2916\ : Odrv12
    port map (
            O => \N__13796\,
            I => charx_if_generate_plus_mult1_un33_sum_i
        );

    \I__2915\ : InMux
    port map (
            O => \N__13793\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_1
        );

    \I__2914\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13786\
        );

    \I__2913\ : InMux
    port map (
            O => \N__13789\,
            I => \N__13783\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__13786\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__13783\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__13778\,
            I => \N__13775\
        );

    \I__2909\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13772\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__13772\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\
        );

    \I__2907\ : InMux
    port map (
            O => \N__13769\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__2906\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13763\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__13763\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\
        );

    \I__2904\ : InMux
    port map (
            O => \N__13760\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__13757\,
            I => \N__13753\
        );

    \I__2902\ : InMux
    port map (
            O => \N__13756\,
            I => \N__13745\
        );

    \I__2901\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13745\
        );

    \I__2900\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13745\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__13745\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0\
        );

    \I__2898\ : InMux
    port map (
            O => \N__13742\,
            I => \N__13739\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__13739\,
            I => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx
        );

    \I__2896\ : InMux
    port map (
            O => \N__13736\,
            I => \N__13733\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__13733\,
            I => \N__13730\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__13730\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\
        );

    \I__2893\ : InMux
    port map (
            O => \N__13727\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__13724\,
            I => \N__13721\
        );

    \I__2891\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13718\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__13718\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0\
        );

    \I__2889\ : InMux
    port map (
            O => \N__13715\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__2888\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13709\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__13709\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\
        );

    \I__2886\ : InMux
    port map (
            O => \N__13706\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__2885\ : InMux
    port map (
            O => \N__13703\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7
        );

    \I__2884\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13697\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__13697\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\
        );

    \I__2882\ : InMux
    port map (
            O => \N__13694\,
            I => \N__13690\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__13693\,
            I => \N__13687\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__13690\,
            I => \N__13679\
        );

    \I__2879\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13675\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__13686\,
            I => \N__13672\
        );

    \I__2877\ : CascadeMux
    port map (
            O => \N__13685\,
            I => \N__13668\
        );

    \I__2876\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13661\
        );

    \I__2875\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13661\
        );

    \I__2874\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13658\
        );

    \I__2873\ : Span4Mux_v
    port map (
            O => \N__13679\,
            I => \N__13655\
        );

    \I__2872\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13652\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__13675\,
            I => \N__13649\
        );

    \I__2870\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13644\
        );

    \I__2869\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13644\
        );

    \I__2868\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13639\
        );

    \I__2867\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13639\
        );

    \I__2866\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13636\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__13661\,
            I => \N__13631\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__13658\,
            I => \N__13631\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__13655\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__13652\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__13649\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__13644\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__13639\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__13636\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2857\ : Odrv12
    port map (
            O => \N__13631\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__13616\,
            I => \N__13610\
        );

    \I__2855\ : InMux
    port map (
            O => \N__13615\,
            I => \N__13606\
        );

    \I__2854\ : InMux
    port map (
            O => \N__13614\,
            I => \N__13602\
        );

    \I__2853\ : InMux
    port map (
            O => \N__13613\,
            I => \N__13599\
        );

    \I__2852\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13596\
        );

    \I__2851\ : InMux
    port map (
            O => \N__13609\,
            I => \N__13593\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__13606\,
            I => \N__13588\
        );

    \I__2849\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13585\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__13602\,
            I => \N__13578\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__13599\,
            I => \N__13578\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__13596\,
            I => \N__13578\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__13593\,
            I => \N__13575\
        );

    \I__2844\ : InMux
    port map (
            O => \N__13592\,
            I => \N__13570\
        );

    \I__2843\ : InMux
    port map (
            O => \N__13591\,
            I => \N__13570\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__13588\,
            I => \N__13565\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__13585\,
            I => \N__13565\
        );

    \I__2840\ : Span4Mux_v
    port map (
            O => \N__13578\,
            I => \N__13562\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__13575\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__13570\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__13565\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__2836\ : Odrv4
    port map (
            O => \N__13562\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__13553\,
            I => \N__13547\
        );

    \I__2834\ : InMux
    port map (
            O => \N__13552\,
            I => \N__13543\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__13551\,
            I => \N__13539\
        );

    \I__2832\ : CascadeMux
    port map (
            O => \N__13550\,
            I => \N__13536\
        );

    \I__2831\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13530\
        );

    \I__2830\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13530\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__13543\,
            I => \N__13527\
        );

    \I__2828\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13524\
        );

    \I__2827\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13517\
        );

    \I__2826\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13517\
        );

    \I__2825\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13517\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__13530\,
            I => \N_520\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__13527\,
            I => \N_520\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__13524\,
            I => \N_520\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__13517\,
            I => \N_520\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__13508\,
            I => \N__13504\
        );

    \I__2819\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13501\
        );

    \I__2818\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13498\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__13501\,
            I => un5_visiblex_i_24
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__13498\,
            I => un5_visiblex_i_24
        );

    \I__2815\ : InMux
    port map (
            O => \N__13493\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_1
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__2813\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13484\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__13484\,
            I => \N__13481\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__13481\,
            I => \column_1_if_generate_plus_mult1_un68_sum_iZ0\
        );

    \I__2810\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__13475\,
            I => if_generate_plus_mult1_un75_sum_cry_2_s
        );

    \I__2808\ : InMux
    port map (
            O => \N__13472\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__2807\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__2805\ : Odrv12
    port map (
            O => \N__13463\,
            I => if_generate_plus_mult1_un68_sum_cry_2_s
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__13460\,
            I => \N__13457\
        );

    \I__2803\ : InMux
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__13454\,
            I => if_generate_plus_mult1_un75_sum_cry_3_s
        );

    \I__2801\ : InMux
    port map (
            O => \N__13451\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__2800\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__13445\,
            I => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\
        );

    \I__2798\ : InMux
    port map (
            O => \N__13442\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__2797\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13436\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2795\ : Odrv12
    port map (
            O => \N__13433\,
            I => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\
        );

    \I__2794\ : InMux
    port map (
            O => \N__13430\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__2793\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13424\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__13424\,
            I => un116_pixel_2_ns_1_2
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__13421\,
            I => \N__13417\
        );

    \I__2790\ : InMux
    port map (
            O => \N__13420\,
            I => \N__13412\
        );

    \I__2789\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13412\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__13412\,
            I => \N__13409\
        );

    \I__2787\ : Odrv12
    port map (
            O => \N__13409\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__2786\ : InMux
    port map (
            O => \N__13406\,
            I => \N__13403\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__13403\,
            I => if_generate_plus_mult1_un75_sum_axb_4_l_fx
        );

    \I__2784\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13397\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__13397\,
            I => \N__13394\
        );

    \I__2782\ : Odrv12
    port map (
            O => \N__13394\,
            I => \beamY_RNII25UDD3_0Z0Z_0\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__13391\,
            I => \un116_pixel_7_ns_1_6_cascade_\
        );

    \I__2780\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13382\
        );

    \I__2779\ : InMux
    port map (
            O => \N__13387\,
            I => \N__13382\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__13382\,
            I => \N__13368\
        );

    \I__2777\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13365\
        );

    \I__2776\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13360\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13360\
        );

    \I__2774\ : InMux
    port map (
            O => \N__13378\,
            I => \N__13353\
        );

    \I__2773\ : InMux
    port map (
            O => \N__13377\,
            I => \N__13353\
        );

    \I__2772\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13353\
        );

    \I__2771\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13350\
        );

    \I__2770\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13343\
        );

    \I__2769\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13343\
        );

    \I__2768\ : InMux
    port map (
            O => \N__13372\,
            I => \N__13343\
        );

    \I__2767\ : InMux
    port map (
            O => \N__13371\,
            I => \N__13340\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__13368\,
            I => font_un3_pixel_29
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__13365\,
            I => font_un3_pixel_29
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__13360\,
            I => font_un3_pixel_29
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__13353\,
            I => font_un3_pixel_29
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__13350\,
            I => font_un3_pixel_29
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__13343\,
            I => font_un3_pixel_29
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__13340\,
            I => font_un3_pixel_29
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__13325\,
            I => \N__13322\
        );

    \I__2758\ : InMux
    port map (
            O => \N__13322\,
            I => \N__13319\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__13319\,
            I => \beamY_RNIBHJ7AMZ0Z_0\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__13316\,
            I => \N__13313\
        );

    \I__2755\ : InMux
    port map (
            O => \N__13313\,
            I => \N__13310\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__13310\,
            I => \N__13307\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__13307\,
            I => \column_1_if_generate_plus_mult1_un75_sum_iZ0\
        );

    \I__2752\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13301\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__13301\,
            I => \G_340\
        );

    \I__2750\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13295\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__13295\,
            I => \G_341\
        );

    \I__2748\ : InMux
    port map (
            O => \N__13292\,
            I => column_1_if_generate_plus_mult1_un82_sum_cry_4
        );

    \I__2747\ : CascadeMux
    port map (
            O => \N__13289\,
            I => \un5_rowlto0_cascade_\
        );

    \I__2746\ : InMux
    port map (
            O => \N__13286\,
            I => \N__13283\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__13283\,
            I => \beamY_RNIJ720T72Z0Z_0\
        );

    \I__2744\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13277\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__13277\,
            I => un116_pixel_5_ns_1_2
        );

    \I__2742\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13271\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__13271\,
            I => \beamY_RNIJDHE4C2Z0Z_1\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__13268\,
            I => \font_un126_pixel_6_am_cascade_\
        );

    \I__2739\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13262\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__13262\,
            I => font_un126_pixel_2_am
        );

    \I__2737\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13256\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__13256\,
            I => \beamX_RNIQ6MATS2Z0Z_0\
        );

    \I__2735\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13250\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__13250\,
            I => \N__13244\
        );

    \I__2733\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13241\
        );

    \I__2732\ : InMux
    port map (
            O => \N__13248\,
            I => \N__13238\
        );

    \I__2731\ : InMux
    port map (
            O => \N__13247\,
            I => \N__13235\
        );

    \I__2730\ : Odrv4
    port map (
            O => \N__13244\,
            I => \un114_pixel_7_1_7__N_11_i_1\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__13241\,
            I => \un114_pixel_7_1_7__N_11_i_1\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__13238\,
            I => \un114_pixel_7_1_7__N_11_i_1\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__13235\,
            I => \un114_pixel_7_1_7__N_11_i_1\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__13226\,
            I => \N_37_cascade_\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__13223\,
            I => \beamY_RNI05CI5A3_1Z0Z_0_cascade_\
        );

    \I__2724\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13217\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__13217\,
            I => \beamY_RNI05CI5A3Z0Z_0\
        );

    \I__2722\ : InMux
    port map (
            O => \N__13214\,
            I => \N__13211\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__13211\,
            I => \beamY_RNII25UDD3_1Z0Z_0\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__13208\,
            I => \un116_pixel_7_ns_1_4_cascade_\
        );

    \I__2719\ : InMux
    port map (
            O => \N__13205\,
            I => \N__13202\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__13202\,
            I => \N__13199\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__13199\,
            I => \beamY_RNIFHEQCT1Z0Z_0\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__13196\,
            I => \beamY_RNIA4V0NM1Z0Z_0_cascade_\
        );

    \I__2715\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13190\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__13190\,
            I => \Pixel_1_r_sn\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__13187\,
            I => \Pixel_1_r_rn_0_cascade_\
        );

    \I__2712\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13181\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__13181\,
            I => \N_396\
        );

    \I__2710\ : IoInMux
    port map (
            O => \N__13178\,
            I => \N__13174\
        );

    \I__2709\ : IoInMux
    port map (
            O => \N__13177\,
            I => \N__13171\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__13174\,
            I => \N__13168\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__13171\,
            I => \N__13165\
        );

    \I__2706\ : Span4Mux_s2_v
    port map (
            O => \N__13168\,
            I => \N__13162\
        );

    \I__2705\ : Span4Mux_s3_v
    port map (
            O => \N__13165\,
            I => \N__13159\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__13162\,
            I => \N__13156\
        );

    \I__2703\ : Span4Mux_h
    port map (
            O => \N__13159\,
            I => \N__13153\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__13156\,
            I => \Pixel_c\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__13153\,
            I => \Pixel_c\
        );

    \I__2700\ : ClkMux
    port map (
            O => \N__13148\,
            I => \N__13103\
        );

    \I__2699\ : ClkMux
    port map (
            O => \N__13147\,
            I => \N__13103\
        );

    \I__2698\ : ClkMux
    port map (
            O => \N__13146\,
            I => \N__13103\
        );

    \I__2697\ : ClkMux
    port map (
            O => \N__13145\,
            I => \N__13103\
        );

    \I__2696\ : ClkMux
    port map (
            O => \N__13144\,
            I => \N__13103\
        );

    \I__2695\ : ClkMux
    port map (
            O => \N__13143\,
            I => \N__13103\
        );

    \I__2694\ : ClkMux
    port map (
            O => \N__13142\,
            I => \N__13103\
        );

    \I__2693\ : ClkMux
    port map (
            O => \N__13141\,
            I => \N__13103\
        );

    \I__2692\ : ClkMux
    port map (
            O => \N__13140\,
            I => \N__13103\
        );

    \I__2691\ : ClkMux
    port map (
            O => \N__13139\,
            I => \N__13103\
        );

    \I__2690\ : ClkMux
    port map (
            O => \N__13138\,
            I => \N__13103\
        );

    \I__2689\ : ClkMux
    port map (
            O => \N__13137\,
            I => \N__13103\
        );

    \I__2688\ : ClkMux
    port map (
            O => \N__13136\,
            I => \N__13103\
        );

    \I__2687\ : ClkMux
    port map (
            O => \N__13135\,
            I => \N__13103\
        );

    \I__2686\ : ClkMux
    port map (
            O => \N__13134\,
            I => \N__13103\
        );

    \I__2685\ : GlobalMux
    port map (
            O => \N__13103\,
            I => \N__13100\
        );

    \I__2684\ : gio2CtrlBuf
    port map (
            O => \N__13100\,
            I => \PixelClock_g\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13094\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__13094\,
            I => \m6Z0Z_1\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13088\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__13088\,
            I => \N__13085\
        );

    \I__2679\ : Span4Mux_h
    port map (
            O => \N__13085\,
            I => \N__13082\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__13082\,
            I => \G_7_0_m2_1\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__13079\,
            I => \beamX_RNI1M3Q1V2Z0Z_0_cascade_\
        );

    \I__2676\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13073\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N_1039_0_0\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__13070\,
            I => \font_un3_pixel_29_cascade_\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__13067\,
            I => \G_7_0_m4_2_1_1_cascade_\
        );

    \I__2672\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13061\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__13061\,
            I => \G_7_0_m4_2_1\
        );

    \I__2670\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13055\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__13055\,
            I => \N__13052\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__13052\,
            I => \beamY_RNINIKJ5A3Z0Z_1\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__13049\,
            I => \beamY_RNI7OTDJ61Z0Z_1_cascade_\
        );

    \I__2666\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13040\
        );

    \I__2665\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13040\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__13040\,
            I => \N__13036\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13039\,
            I => \N__13033\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__13036\,
            I => un4_row
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__13033\,
            I => un4_row
        );

    \I__2660\ : InMux
    port map (
            O => \N__13028\,
            I => \N__13025\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__13025\,
            I => \N__13022\
        );

    \I__2658\ : Span4Mux_h
    port map (
            O => \N__13022\,
            I => \N__13019\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__13019\,
            I => \beamY_RNIPG1SS93Z0Z_2\
        );

    \I__2656\ : InMux
    port map (
            O => \N__13016\,
            I => \N__13013\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__13013\,
            I => \N_23_0\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13010\,
            I => \N__13007\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__13007\,
            I => \N_15_0\
        );

    \I__2652\ : InMux
    port map (
            O => \N__13004\,
            I => \N__13001\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13001\,
            I => \N_342_0_0\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__12998\,
            I => \N_1045_0_cascade_\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__12995\,
            I => \N__12992\
        );

    \I__2648\ : InMux
    port map (
            O => \N__12992\,
            I => \N__12989\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__12989\,
            I => \column_1_if_generate_plus_mult1_un61_sum_iZ0\
        );

    \I__2646\ : InMux
    port map (
            O => \N__12986\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__12983\,
            I => \N__12980\
        );

    \I__2644\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12977\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__12977\,
            I => \N__12974\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__12974\,
            I => \N__12971\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__12971\,
            I => if_generate_plus_mult1_un61_sum_cry_2_s
        );

    \I__2640\ : InMux
    port map (
            O => \N__12968\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__2639\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12959\
        );

    \I__2638\ : InMux
    port map (
            O => \N__12964\,
            I => \N__12959\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__12959\,
            I => un5_rowlto3_i
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__12956\,
            I => \N__12953\
        );

    \I__2635\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12950\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__12950\,
            I => \N__12947\
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__12947\,
            I => if_generate_plus_mult1_un61_sum_cry_3_s
        );

    \I__2632\ : InMux
    port map (
            O => \N__12944\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__2631\ : InMux
    port map (
            O => \N__12941\,
            I => \N__12938\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__12938\,
            I => \N__12935\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__12935\,
            I => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\
        );

    \I__2628\ : InMux
    port map (
            O => \N__12932\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__2627\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12926\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__12926\,
            I => \Pixel_3_sqmuxa\
        );

    \I__2625\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12920\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__12920\,
            I => \un114_pixel_6_1_5__font_un126_pixel_m_4\
        );

    \I__2623\ : CascadeMux
    port map (
            O => \N__12917\,
            I => \N__12914\
        );

    \I__2622\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12911\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__2620\ : Span4Mux_h
    port map (
            O => \N__12908\,
            I => \N__12905\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__12905\,
            I => un1_beamy_0_0
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__12902\,
            I => \un116_pixel_5_amZ0Z_6_cascade_\
        );

    \I__2617\ : InMux
    port map (
            O => \N__12899\,
            I => \N__12896\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__12896\,
            I => \un116_pixel_5_bmZ0Z_6\
        );

    \I__2615\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12889\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__12892\,
            I => \N__12886\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__12889\,
            I => \N__12883\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12880\
        );

    \I__2611\ : Span4Mux_h
    port map (
            O => \N__12883\,
            I => \N__12877\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__12880\,
            I => un15_beamy
        );

    \I__2609\ : Odrv4
    port map (
            O => \N__12877\,
            I => un15_beamy
        );

    \I__2608\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12869\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__12869\,
            I => \N__12866\
        );

    \I__2606\ : Span4Mux_v
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__12863\,
            I => \un114_pixel_6_1_5__g0Z0Z_0\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__12860\,
            I => \un114_pixel_6_1_5__font_un126_pixel_mZ0Z_1_cascade_\
        );

    \I__2603\ : InMux
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__12854\,
            I => \N__12851\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__12851\,
            I => \N__12848\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__12848\,
            I => \un114_pixel_6_1_5__font_un126_pixel_m_4_1_0\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__12845\,
            I => \un114_pixel_6_1_5__g0_2Z0Z_0_cascade_\
        );

    \I__2598\ : InMux
    port map (
            O => \N__12842\,
            I => \N__12839\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__12839\,
            I => \N__12836\
        );

    \I__2596\ : Span4Mux_v
    port map (
            O => \N__12836\,
            I => \N__12833\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__12833\,
            I => \un114_pixel_6_1_5__font_un126_pixel_m_4_1_1_0\
        );

    \I__2594\ : InMux
    port map (
            O => \N__12830\,
            I => \N__12827\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__12827\,
            I => \N__12824\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__12824\,
            I => \N__12821\
        );

    \I__2591\ : Odrv4
    port map (
            O => \N__12821\,
            I => \un114_pixel_6_1_5__g0_1_0\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__12818\,
            I => \un114_pixel_6_1_5__g1Z0Z_0_cascade_\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__12815\,
            I => \N__12812\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12809\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__12809\,
            I => charx_if_generate_plus_mult1_un26_sum_s_2_sf
        );

    \I__2586\ : InMux
    port map (
            O => \N__12806\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_1
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__2584\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12797\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__12797\,
            I => \un5_visiblex_cry_8_c_RNI1D62Z0Z_2\
        );

    \I__2582\ : InMux
    port map (
            O => \N__12794\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__2581\ : InMux
    port map (
            O => \N__12791\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_3
        );

    \I__2580\ : InMux
    port map (
            O => \N__12788\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_4
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__12785\,
            I => \N__12782\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12779\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__12779\,
            I => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__2575\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__12770\,
            I => un5_visiblex_i_25
        );

    \I__2573\ : InMux
    port map (
            O => \N__12767\,
            I => \N__12762\
        );

    \I__2572\ : InMux
    port map (
            O => \N__12766\,
            I => \N__12759\
        );

    \I__2571\ : InMux
    port map (
            O => \N__12765\,
            I => \N__12756\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__12762\,
            I => column_1_if_generate_plus_mult1_un47_sum0_5
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__12759\,
            I => column_1_if_generate_plus_mult1_un47_sum0_5
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__12756\,
            I => column_1_if_generate_plus_mult1_un47_sum0_5
        );

    \I__2567\ : CascadeMux
    port map (
            O => \N__12749\,
            I => \N__12745\
        );

    \I__2566\ : CascadeMux
    port map (
            O => \N__12748\,
            I => \N__12742\
        );

    \I__2565\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12739\
        );

    \I__2564\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12736\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__12739\,
            I => column_1_if_generate_plus_mult1_un47_sum1_5
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__12736\,
            I => column_1_if_generate_plus_mult1_un47_sum1_5
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__12731\,
            I => \N__12728\
        );

    \I__2560\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12725\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__12725\,
            I => \un114_pixel_6_1_5__un4_rowZ0Z_0\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__2557\ : InMux
    port map (
            O => \N__12719\,
            I => \N__12716\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__12716\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i
        );

    \I__2555\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12710\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__12710\,
            I => \N__12707\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__12707\,
            I => column_1_if_generate_plus_mult1_un47_sum0_2
        );

    \I__2552\ : InMux
    port map (
            O => \N__12704\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_1
        );

    \I__2551\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12698\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__12698\,
            I => column_1_if_generate_plus_mult1_un47_sum0_3
        );

    \I__2549\ : InMux
    port map (
            O => \N__12695\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_2
        );

    \I__2548\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12689\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__12689\,
            I => column_1_if_generate_plus_mult1_un47_sum0_4
        );

    \I__2546\ : InMux
    port map (
            O => \N__12686\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_3
        );

    \I__2545\ : InMux
    port map (
            O => \N__12683\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_4
        );

    \I__2544\ : InMux
    port map (
            O => \N__12680\,
            I => \N__12677\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__12677\,
            I => if_generate_plus_mult1_un47_sum_0_cry_3_ma
        );

    \I__2542\ : InMux
    port map (
            O => \N__12674\,
            I => \N__12671\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__12671\,
            I => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2539\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__12662\,
            I => \N_200_0_i\
        );

    \I__2537\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__12656\,
            I => \un116_pixel_4_bmZ0Z_1\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__12653\,
            I => \un116_pixel_4_amZ0Z_1_cascade_\
        );

    \I__2534\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12647\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__12647\,
            I => un116_pixel_3_ns_1_1
        );

    \I__2532\ : InMux
    port map (
            O => \N__12644\,
            I => \N__12641\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__12641\,
            I => \N__12638\
        );

    \I__2530\ : Odrv12
    port map (
            O => \N__12638\,
            I => \beamY_RNIHIRVUS1Z0Z_1\
        );

    \I__2529\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12632\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__12632\,
            I => \un116_pixel_1_bmZ0Z_1\
        );

    \I__2527\ : InMux
    port map (
            O => \N__12629\,
            I => \N__12626\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__12626\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421\
        );

    \I__2525\ : InMux
    port map (
            O => \N__12623\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__12620\,
            I => \N__12617\
        );

    \I__2523\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12614\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__12614\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1\
        );

    \I__2521\ : InMux
    port map (
            O => \N__12611\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__2520\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12605\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__12605\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8
        );

    \I__2518\ : InMux
    port map (
            O => \N__12602\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__2517\ : InMux
    port map (
            O => \N__12599\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__12596\,
            I => \N__12592\
        );

    \I__2515\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12588\
        );

    \I__2514\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12583\
        );

    \I__2513\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12583\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__12588\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__12583\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\
        );

    \I__2510\ : InMux
    port map (
            O => \N__12578\,
            I => \N__12572\
        );

    \I__2509\ : InMux
    port map (
            O => \N__12577\,
            I => \N__12572\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__12572\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__12569\,
            I => \un114_pixel_3_i_a3_7_cascade_\
        );

    \I__2506\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__12563\,
            I => \N__12559\
        );

    \I__2504\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12556\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__12559\,
            I => column_0001_0
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__12556\,
            I => column_0001_0
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__12551\,
            I => \un116_pixel_3_ns_1_2_cascade_\
        );

    \I__2500\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__12545\,
            I => \beamY_RNIDVSK5A3Z0Z_1\
        );

    \I__2498\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12539\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__12539\,
            I => \N_13_0\
        );

    \I__2496\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12533\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__2494\ : Odrv4
    port map (
            O => \N__12530\,
            I => \un114_pixel_0_1__N_6_mux_0\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__12527\,
            I => \un116_pixel_1_amZ0Z_1_cascade_\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__12524\,
            I => \un116_pixel_3_bmZ0Z_6_cascade_\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__12521\,
            I => \beamY_RNISJITRQ2Z0Z_1_cascade_\
        );

    \I__2490\ : InMux
    port map (
            O => \N__12518\,
            I => \N__12515\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12515\,
            I => \N_12_0\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__12512\,
            I => \N_248_0_cascade_\
        );

    \I__2487\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__12506\,
            I => un116_pixel_3_ns_1_0_6
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \N__12500\
        );

    \I__2484\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12497\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__12497\,
            I => \N_25_mux\
        );

    \I__2482\ : InMux
    port map (
            O => \N__12494\,
            I => \N__12491\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__12491\,
            I => \N__12488\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__12488\,
            I => \N__12485\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__12485\,
            I => font_un28_pixel_0_0_29
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__12482\,
            I => \un114_pixel_6_1_5__un116_pixel_3_1_0_0_7_cascade_\
        );

    \I__2477\ : InMux
    port map (
            O => \N__12479\,
            I => \N__12476\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__12476\,
            I => \N_14_0\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__12473\,
            I => \column_0111_0_cascade_\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__12470\,
            I => \beamY_RNI05CI5A3_0Z0Z_0_cascade_\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__12467\,
            I => \beamY_RNIBABJS01Z0Z_1_cascade_\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__12464\,
            I => \N_21_0_cascade_\
        );

    \I__2471\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__12458\,
            I => \N_22_0\
        );

    \I__2469\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12452\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__12452\,
            I => column_0111_0
        );

    \I__2467\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12446\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__12446\,
            I => \N__12443\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__12443\,
            I => chessboardpixel_un174_pixel_0_1
        );

    \I__2464\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12437\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__12437\,
            I => chessboardpixel_un200_pixel_0_1
        );

    \I__2462\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__12431\,
            I => \un114_pixel_6_1_5__un4_row_7Z0Z_1\
        );

    \I__2460\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12425\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__12425\,
            I => \N_357_0\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__12422\,
            I => \N_18_0_cascade_\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__12419\,
            I => \N_7_0_cascade_\
        );

    \I__2456\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12410\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__12410\,
            I => if_generate_plus_mult1_un54_sum_axb_4_l_fx
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__2452\ : InMux
    port map (
            O => \N__12404\,
            I => \N__12400\
        );

    \I__2451\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12397\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__12400\,
            I => \N__12391\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__12397\,
            I => \N__12391\
        );

    \I__2448\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12388\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__12391\,
            I => \N_571_i\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__12388\,
            I => \N_571_i\
        );

    \I__2445\ : InMux
    port map (
            O => \N__12383\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__2444\ : InMux
    port map (
            O => \N__12380\,
            I => \N__12377\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__12377\,
            I => \N__12374\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__12374\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\
        );

    \I__2441\ : InMux
    port map (
            O => \N__12371\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__12368\,
            I => \if_generate_plus_mult1_un54_sum_s_5_cascade_\
        );

    \I__2439\ : InMux
    port map (
            O => \N__12365\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__2438\ : InMux
    port map (
            O => \N__12362\,
            I => \N__12357\
        );

    \I__2437\ : InMux
    port map (
            O => \N__12361\,
            I => \N__12354\
        );

    \I__2436\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12351\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__12357\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__12354\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__12351\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__12344\,
            I => \N__12341\
        );

    \I__2431\ : InMux
    port map (
            O => \N__12341\,
            I => \N__12338\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__12338\,
            I => if_generate_plus_mult1_un54_sum_cry_2_s
        );

    \I__2429\ : InMux
    port map (
            O => \N__12335\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__2428\ : InMux
    port map (
            O => \N__12332\,
            I => \N__12326\
        );

    \I__2427\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12326\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__12326\,
            I => column_1_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__12323\,
            I => \N__12320\
        );

    \I__2424\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12317\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__12317\,
            I => if_generate_plus_mult1_un54_sum_cry_3_s
        );

    \I__2422\ : InMux
    port map (
            O => \N__12314\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__2421\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12308\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__12308\,
            I => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\
        );

    \I__2419\ : InMux
    port map (
            O => \N__12305\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__12302\,
            I => \N__12299\
        );

    \I__2417\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12296\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__12296\,
            I => \N_562_i\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__12293\,
            I => \N__12290\
        );

    \I__2414\ : InMux
    port map (
            O => \N__12290\,
            I => \N__12287\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__12287\,
            I => \N_11_0_i\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__12284\,
            I => \N__12281\
        );

    \I__2411\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12278\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__12278\,
            I => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx
        );

    \I__2409\ : InMux
    port map (
            O => \N__12275\,
            I => \N__12272\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12267\
        );

    \I__2407\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12264\
        );

    \I__2406\ : InMux
    port map (
            O => \N__12270\,
            I => \N__12261\
        );

    \I__2405\ : Span4Mux_h
    port map (
            O => \N__12267\,
            I => \N__12251\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__12264\,
            I => \N__12248\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__12261\,
            I => \N__12245\
        );

    \I__2402\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12237\
        );

    \I__2401\ : InMux
    port map (
            O => \N__12259\,
            I => \N__12237\
        );

    \I__2400\ : InMux
    port map (
            O => \N__12258\,
            I => \N__12237\
        );

    \I__2399\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12230\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12256\,
            I => \N__12227\
        );

    \I__2397\ : InMux
    port map (
            O => \N__12255\,
            I => \N__12224\
        );

    \I__2396\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12221\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__12251\,
            I => \N__12216\
        );

    \I__2394\ : Span4Mux_h
    port map (
            O => \N__12248\,
            I => \N__12216\
        );

    \I__2393\ : Span4Mux_v
    port map (
            O => \N__12245\,
            I => \N__12213\
        );

    \I__2392\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12210\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__12237\,
            I => \N__12207\
        );

    \I__2390\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12198\
        );

    \I__2389\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12198\
        );

    \I__2388\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12198\
        );

    \I__2387\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12198\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__12230\,
            I => \N__12191\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__12227\,
            I => \N__12191\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__12224\,
            I => \N__12191\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__12221\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__12216\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__12213\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__12210\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__12207\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__12198\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2377\ : Odrv12
    port map (
            O => \N__12191\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2376\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12170\
        );

    \I__2375\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12165\
        );

    \I__2374\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12162\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__12173\,
            I => \N__12159\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__12170\,
            I => \N__12155\
        );

    \I__2371\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12151\
        );

    \I__2370\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12148\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__12165\,
            I => \N__12143\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__12162\,
            I => \N__12143\
        );

    \I__2367\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12138\
        );

    \I__2366\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12138\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__12155\,
            I => \N__12135\
        );

    \I__2364\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12132\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__12151\,
            I => \N__12129\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__12148\,
            I => \N__12126\
        );

    \I__2361\ : Odrv12
    port map (
            O => \N__12143\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12138\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__12135\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__12132\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__12129\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__12126\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3
        );

    \I__2355\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12109\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__12112\,
            I => \N__12105\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__12109\,
            I => \N__12098\
        );

    \I__2352\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12095\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12092\
        );

    \I__2350\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12085\
        );

    \I__2349\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12085\
        );

    \I__2348\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12077\
        );

    \I__2347\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12077\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__12098\,
            I => \N__12074\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__12095\,
            I => \N__12071\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__12092\,
            I => \N__12068\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12063\
        );

    \I__2342\ : InMux
    port map (
            O => \N__12090\,
            I => \N__12063\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__12085\,
            I => \N__12055\
        );

    \I__2340\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12050\
        );

    \I__2339\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12050\
        );

    \I__2338\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12047\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__12077\,
            I => \N__12044\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__12074\,
            I => \N__12041\
        );

    \I__2335\ : Span4Mux_v
    port map (
            O => \N__12071\,
            I => \N__12034\
        );

    \I__2334\ : Span4Mux_v
    port map (
            O => \N__12068\,
            I => \N__12034\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__12063\,
            I => \N__12034\
        );

    \I__2332\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12027\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12061\,
            I => \N__12027\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12027\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12022\
        );

    \I__2328\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12022\
        );

    \I__2327\ : Span4Mux_h
    port map (
            O => \N__12055\,
            I => \N__12019\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__12050\,
            I => \N__12012\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__12047\,
            I => \N__12012\
        );

    \I__2324\ : Span12Mux_s2_v
    port map (
            O => \N__12044\,
            I => \N__12012\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__12041\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__12034\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__12027\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__12022\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__12019\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2318\ : Odrv12
    port map (
            O => \N__12012\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__11999\,
            I => \N__11996\
        );

    \I__2316\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11993\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__11993\,
            I => \un114_pixel_6_1_5__un4_rowZ0Z_2\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__11990\,
            I => \N__11987\
        );

    \I__2313\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11984\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__11984\,
            I => if_generate_plus_mult1_un47_sum_m_1
        );

    \I__2311\ : InMux
    port map (
            O => \N__11981\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__2310\ : InMux
    port map (
            O => \N__11978\,
            I => \N__11975\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__11975\,
            I => \N__11971\
        );

    \I__2308\ : InMux
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__11971\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__11968\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__11963\,
            I => \N__11960\
        );

    \I__2304\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__11957\,
            I => \N__11954\
        );

    \I__2302\ : Odrv12
    port map (
            O => \N__11954\,
            I => if_generate_plus_mult1_un47_sum_m_2
        );

    \I__2301\ : InMux
    port map (
            O => \N__11951\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__2300\ : InMux
    port map (
            O => \N__11948\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_4
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__11945\,
            I => \column_1_if_generate_plus_mult1_un47_sum1_5_cascade_\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__11942\,
            I => \N__11939\
        );

    \I__2297\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__11936\,
            I => un5_visiblex_i_0_25
        );

    \I__2295\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11930\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__11930\,
            I => charx_if_generate_plus_mult1_un26_sum_axb_3_i
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__11927\,
            I => \N__11924\
        );

    \I__2292\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11921\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__2290\ : Odrv4
    port map (
            O => \N__11918\,
            I => column_1_if_generate_plus_mult1_un47_sum1_4
        );

    \I__2289\ : InMux
    port map (
            O => \N__11915\,
            I => \N__11912\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__11912\,
            I => column_1_if_generate_plus_mult1_un47_sum1_3
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__11909\,
            I => \if_generate_plus_mult1_un47_sum_m_5_cascade_\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__11906\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__11903\,
            I => \N__11900\
        );

    \I__2284\ : InMux
    port map (
            O => \N__11900\,
            I => \N__11897\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__11897\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2\
        );

    \I__2282\ : InMux
    port map (
            O => \N__11894\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__2281\ : InMux
    port map (
            O => \N__11891\,
            I => \N__11888\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__11888\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__2279\ : InMux
    port map (
            O => \N__11885\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__2278\ : InMux
    port map (
            O => \N__11882\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__2277\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11874\
        );

    \I__2276\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11869\
        );

    \I__2275\ : InMux
    port map (
            O => \N__11877\,
            I => \N__11869\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__11874\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__11869\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__11864\,
            I => \N__11861\
        );

    \I__2271\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11858\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__11858\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i
        );

    \I__2269\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11849\
        );

    \I__2268\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11849\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__11849\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__2266\ : InMux
    port map (
            O => \N__11846\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_1
        );

    \I__2265\ : InMux
    port map (
            O => \N__11843\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_2
        );

    \I__2264\ : InMux
    port map (
            O => \N__11840\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_3
        );

    \I__2263\ : InMux
    port map (
            O => \N__11837\,
            I => \N__11834\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__11834\,
            I => g1_0_1
        );

    \I__2261\ : CascadeMux
    port map (
            O => \N__11831\,
            I => \N__11824\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__11830\,
            I => \N__11819\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__11829\,
            I => \N__11816\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__11828\,
            I => \N__11812\
        );

    \I__2257\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11805\
        );

    \I__2256\ : InMux
    port map (
            O => \N__11824\,
            I => \N__11800\
        );

    \I__2255\ : InMux
    port map (
            O => \N__11823\,
            I => \N__11800\
        );

    \I__2254\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11797\
        );

    \I__2253\ : InMux
    port map (
            O => \N__11819\,
            I => \N__11789\
        );

    \I__2252\ : InMux
    port map (
            O => \N__11816\,
            I => \N__11789\
        );

    \I__2251\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11786\
        );

    \I__2250\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11783\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__11811\,
            I => \N__11777\
        );

    \I__2248\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11773\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__11809\,
            I => \N__11769\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11766\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__11805\,
            I => \N__11759\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__11800\,
            I => \N__11759\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__11797\,
            I => \N__11759\
        );

    \I__2242\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11756\
        );

    \I__2241\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11751\
        );

    \I__2240\ : InMux
    port map (
            O => \N__11794\,
            I => \N__11751\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__11789\,
            I => \N__11748\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__11786\,
            I => \N__11743\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__11783\,
            I => \N__11743\
        );

    \I__2236\ : InMux
    port map (
            O => \N__11782\,
            I => \N__11740\
        );

    \I__2235\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11737\
        );

    \I__2234\ : InMux
    port map (
            O => \N__11780\,
            I => \N__11734\
        );

    \I__2233\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11729\
        );

    \I__2232\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11729\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__11773\,
            I => \N__11726\
        );

    \I__2230\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11721\
        );

    \I__2229\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11721\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__11766\,
            I => \N__11718\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__11759\,
            I => \N__11715\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__11756\,
            I => \N__11698\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__11751\,
            I => \N__11698\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__11748\,
            I => \N__11698\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__11743\,
            I => \N__11698\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__11740\,
            I => \N__11698\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__11737\,
            I => \N__11698\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__11734\,
            I => \N__11698\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__11729\,
            I => \N__11698\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__11726\,
            I => \N__11693\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__11721\,
            I => \N__11693\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__11718\,
            I => \N__11686\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__11715\,
            I => \N__11686\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__11698\,
            I => \N__11686\
        );

    \I__2213\ : Span4Mux_h
    port map (
            O => \N__11693\,
            I => \N__11683\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__11686\,
            I => \beamYZ0Z_3\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__11683\,
            I => \beamYZ0Z_3\
        );

    \I__2210\ : InMux
    port map (
            O => \N__11678\,
            I => \N__11674\
        );

    \I__2209\ : InMux
    port map (
            O => \N__11677\,
            I => \N__11668\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__11674\,
            I => \N__11665\
        );

    \I__2207\ : InMux
    port map (
            O => \N__11673\,
            I => \N__11660\
        );

    \I__2206\ : InMux
    port map (
            O => \N__11672\,
            I => \N__11660\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__11671\,
            I => \N__11654\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__11668\,
            I => \N__11650\
        );

    \I__2203\ : Span4Mux_h
    port map (
            O => \N__11665\,
            I => \N__11645\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__11660\,
            I => \N__11645\
        );

    \I__2201\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11642\
        );

    \I__2200\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11633\
        );

    \I__2199\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11633\
        );

    \I__2198\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11633\
        );

    \I__2197\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11633\
        );

    \I__2196\ : Span12Mux_s4_v
    port map (
            O => \N__11650\,
            I => \N__11630\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__11645\,
            I => \N__11627\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__11642\,
            I => \N__11622\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__11633\,
            I => \N__11622\
        );

    \I__2192\ : Odrv12
    port map (
            O => \N__11630\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__11627\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2190\ : Odrv12
    port map (
            O => \N__11622\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i
        );

    \I__2189\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__11612\,
            I => g2
        );

    \I__2187\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__11606\,
            I => m511_0_o2_1
        );

    \I__2185\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11597\
        );

    \I__2184\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11597\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__11597\,
            I => \N__11594\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__11594\,
            I => \N__11585\
        );

    \I__2181\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11582\
        );

    \I__2180\ : InMux
    port map (
            O => \N__11592\,
            I => \N__11579\
        );

    \I__2179\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11570\
        );

    \I__2178\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11570\
        );

    \I__2177\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11570\
        );

    \I__2176\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11570\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__11585\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__11582\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__11579\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__11570\,
            I => chary_if_generate_plus_mult1_un68_sum_axbxc5_0
        );

    \I__2171\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11558\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__11558\,
            I => \N_80_i\
        );

    \I__2169\ : CEMux
    port map (
            O => \N__11555\,
            I => \N__11550\
        );

    \I__2168\ : CEMux
    port map (
            O => \N__11554\,
            I => \N__11547\
        );

    \I__2167\ : InMux
    port map (
            O => \N__11553\,
            I => \N__11539\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__11550\,
            I => \N__11534\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__11547\,
            I => \N__11534\
        );

    \I__2164\ : CEMux
    port map (
            O => \N__11546\,
            I => \N__11531\
        );

    \I__2163\ : CEMux
    port map (
            O => \N__11545\,
            I => \N__11527\
        );

    \I__2162\ : CEMux
    port map (
            O => \N__11544\,
            I => \N__11524\
        );

    \I__2161\ : CEMux
    port map (
            O => \N__11543\,
            I => \N__11521\
        );

    \I__2160\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11518\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__11539\,
            I => \N__11515\
        );

    \I__2158\ : Span4Mux_v
    port map (
            O => \N__11534\,
            I => \N__11510\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__11531\,
            I => \N__11510\
        );

    \I__2156\ : CEMux
    port map (
            O => \N__11530\,
            I => \N__11504\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__11527\,
            I => \N__11501\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__11524\,
            I => \N__11496\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__11521\,
            I => \N__11496\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__11518\,
            I => \N__11491\
        );

    \I__2151\ : Span4Mux_v
    port map (
            O => \N__11515\,
            I => \N__11491\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__11510\,
            I => \N__11488\
        );

    \I__2149\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11485\
        );

    \I__2148\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11482\
        );

    \I__2147\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11479\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__11504\,
            I => \N__11476\
        );

    \I__2145\ : Span12Mux_s6_v
    port map (
            O => \N__11501\,
            I => \N__11473\
        );

    \I__2144\ : Span4Mux_v
    port map (
            O => \N__11496\,
            I => \N__11466\
        );

    \I__2143\ : Span4Mux_v
    port map (
            O => \N__11491\,
            I => \N__11466\
        );

    \I__2142\ : Span4Mux_v
    port map (
            O => \N__11488\,
            I => \N__11466\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__11485\,
            I => un3_beamx_0
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__11482\,
            I => un3_beamx_0
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__11479\,
            I => un3_beamx_0
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__11476\,
            I => un3_beamx_0
        );

    \I__2137\ : Odrv12
    port map (
            O => \N__11473\,
            I => un3_beamx_0
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__11466\,
            I => un3_beamx_0
        );

    \I__2135\ : InMux
    port map (
            O => \N__11453\,
            I => \N__11450\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__11450\,
            I => \N__11443\
        );

    \I__2133\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11440\
        );

    \I__2132\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11437\
        );

    \I__2131\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11434\
        );

    \I__2130\ : InMux
    port map (
            O => \N__11446\,
            I => \N__11431\
        );

    \I__2129\ : Span12Mux_s3_h
    port map (
            O => \N__11443\,
            I => \N__11422\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__11440\,
            I => \N__11422\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__11437\,
            I => \N__11419\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__11434\,
            I => \N__11416\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__11431\,
            I => \N__11413\
        );

    \I__2124\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11404\
        );

    \I__2123\ : InMux
    port map (
            O => \N__11429\,
            I => \N__11404\
        );

    \I__2122\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11404\
        );

    \I__2121\ : InMux
    port map (
            O => \N__11427\,
            I => \N__11404\
        );

    \I__2120\ : Span12Mux_s8_h
    port map (
            O => \N__11422\,
            I => \N__11401\
        );

    \I__2119\ : Span4Mux_h
    port map (
            O => \N__11419\,
            I => \N__11396\
        );

    \I__2118\ : Span4Mux_s3_h
    port map (
            O => \N__11416\,
            I => \N__11396\
        );

    \I__2117\ : Span4Mux_s3_h
    port map (
            O => \N__11413\,
            I => \N__11393\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__11404\,
            I => \N__11390\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__11401\,
            I => un5_beamx_0
        );

    \I__2114\ : Odrv4
    port map (
            O => \N__11396\,
            I => un5_beamx_0
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__11393\,
            I => un5_beamx_0
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__11390\,
            I => un5_beamx_0
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__11381\,
            I => \N__11371\
        );

    \I__2110\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11362\
        );

    \I__2109\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11359\
        );

    \I__2108\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11356\
        );

    \I__2107\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11353\
        );

    \I__2106\ : InMux
    port map (
            O => \N__11376\,
            I => \N__11348\
        );

    \I__2105\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11348\
        );

    \I__2104\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11345\
        );

    \I__2103\ : InMux
    port map (
            O => \N__11371\,
            I => \N__11342\
        );

    \I__2102\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11337\
        );

    \I__2101\ : InMux
    port map (
            O => \N__11369\,
            I => \N__11337\
        );

    \I__2100\ : InMux
    port map (
            O => \N__11368\,
            I => \N__11334\
        );

    \I__2099\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11325\
        );

    \I__2098\ : InMux
    port map (
            O => \N__11366\,
            I => \N__11322\
        );

    \I__2097\ : InMux
    port map (
            O => \N__11365\,
            I => \N__11318\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__11362\,
            I => \N__11315\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__11359\,
            I => \N__11312\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__11356\,
            I => \N__11307\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__11353\,
            I => \N__11307\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__11348\,
            I => \N__11304\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__11345\,
            I => \N__11295\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11295\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__11337\,
            I => \N__11295\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__11334\,
            I => \N__11295\
        );

    \I__2087\ : InMux
    port map (
            O => \N__11333\,
            I => \N__11288\
        );

    \I__2086\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11288\
        );

    \I__2085\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11288\
        );

    \I__2084\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11285\
        );

    \I__2083\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11280\
        );

    \I__2082\ : InMux
    port map (
            O => \N__11328\,
            I => \N__11280\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__11325\,
            I => \N__11277\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__11322\,
            I => \N__11274\
        );

    \I__2079\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11271\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__11318\,
            I => \N__11268\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__11315\,
            I => \N__11255\
        );

    \I__2076\ : Span4Mux_v
    port map (
            O => \N__11312\,
            I => \N__11255\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__11307\,
            I => \N__11255\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__11304\,
            I => \N__11255\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__11295\,
            I => \N__11255\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__11288\,
            I => \N__11255\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__11285\,
            I => \N__11250\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__11280\,
            I => \N__11250\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__11277\,
            I => \N__11245\
        );

    \I__2068\ : Span4Mux_v
    port map (
            O => \N__11274\,
            I => \N__11245\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__11271\,
            I => \N__11242\
        );

    \I__2066\ : Span4Mux_h
    port map (
            O => \N__11268\,
            I => \N__11237\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__11255\,
            I => \N__11237\
        );

    \I__2064\ : Span4Mux_h
    port map (
            O => \N__11250\,
            I => \N__11234\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__11245\,
            I => \beamYZ0Z_2\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__11242\,
            I => \beamYZ0Z_2\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__11237\,
            I => \beamYZ0Z_2\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__11234\,
            I => \beamYZ0Z_2\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11225\,
            I => \N__11222\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__11222\,
            I => \N__11219\
        );

    \I__2057\ : Odrv12
    port map (
            O => \N__11219\,
            I => chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_0
        );

    \I__2056\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11212\
        );

    \I__2055\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11209\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__11212\,
            I => \beamY_RNIJH2N2PZ0Z_3\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__11209\,
            I => \beamY_RNIJH2N2PZ0Z_3\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__2051\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11198\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__11198\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1\
        );

    \I__2049\ : InMux
    port map (
            O => \N__11195\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2048\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11185\
        );

    \I__2047\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11185\
        );

    \I__2046\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11182\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__11185\,
            I => \N__11179\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__11182\,
            I => un1_beamx_2
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__11179\,
            I => un1_beamx_2
        );

    \I__2042\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11163\
        );

    \I__2041\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11163\
        );

    \I__2040\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11163\
        );

    \I__2039\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11159\
        );

    \I__2038\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11156\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__11163\,
            I => \N__11153\
        );

    \I__2036\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11150\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__11159\,
            I => \beamXZ0Z_7\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__11156\,
            I => \beamXZ0Z_7\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__11153\,
            I => \beamXZ0Z_7\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__11150\,
            I => \beamXZ0Z_7\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__11141\,
            I => \N__11135\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__11140\,
            I => \N__11132\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__11139\,
            I => \N__11129\
        );

    \I__2028\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11126\
        );

    \I__2027\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11123\
        );

    \I__2026\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11120\
        );

    \I__2025\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11117\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__11126\,
            I => \beamXZ0Z_10\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__11123\,
            I => \beamXZ0Z_10\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__11120\,
            I => \beamXZ0Z_10\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__11117\,
            I => \beamXZ0Z_10\
        );

    \I__2020\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__11105\,
            I => un1_beamxlt10_0
        );

    \I__2018\ : IoInMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__11099\,
            I => \N__11095\
        );

    \I__2016\ : IoInMux
    port map (
            O => \N__11098\,
            I => \N__11092\
        );

    \I__2015\ : Span4Mux_s1_v
    port map (
            O => \N__11095\,
            I => \N__11089\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__11092\,
            I => \N__11086\
        );

    \I__2013\ : Sp12to4
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__2012\ : Span4Mux_s3_v
    port map (
            O => \N__11086\,
            I => \N__11080\
        );

    \I__2011\ : Span12Mux_s6_h
    port map (
            O => \N__11083\,
            I => \N__11077\
        );

    \I__2010\ : Span4Mux_v
    port map (
            O => \N__11080\,
            I => \N__11074\
        );

    \I__2009\ : Odrv12
    port map (
            O => \N__11077\,
            I => \HSync_c\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__11074\,
            I => \HSync_c\
        );

    \I__2007\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__11063\,
            I => \un114_pixel_6_1_5__un4_rowZ0Z_5\
        );

    \I__2004\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11056\
        );

    \I__2003\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11053\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__11056\,
            I => \N__11044\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__11053\,
            I => \N__11044\
        );

    \I__2000\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11035\
        );

    \I__1999\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11035\
        );

    \I__1998\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11035\
        );

    \I__1997\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11035\
        );

    \I__1996\ : Span4Mux_v
    port map (
            O => \N__11044\,
            I => \N__11032\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__11035\,
            I => \N__11029\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__11032\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__11029\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__11024\,
            I => \N__11021\
        );

    \I__1991\ : InMux
    port map (
            O => \N__11021\,
            I => \N__11018\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__11018\,
            I => \N__11014\
        );

    \I__1989\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11011\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__11014\,
            I => \N__11005\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__11011\,
            I => \N__11002\
        );

    \I__1986\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10997\
        );

    \I__1985\ : InMux
    port map (
            O => \N__11009\,
            I => \N__10997\
        );

    \I__1984\ : InMux
    port map (
            O => \N__11008\,
            I => \N__10994\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__11005\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__11002\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__10997\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__10994\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\
        );

    \I__1979\ : InMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__10982\,
            I => \N__10979\
        );

    \I__1977\ : Span4Mux_h
    port map (
            O => \N__10979\,
            I => \N__10976\
        );

    \I__1976\ : Odrv4
    port map (
            O => \N__10976\,
            I => if_generate_plus_mult1_un75_sum_axbxc5
        );

    \I__1975\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10970\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__10970\,
            I => \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_3\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__10967\,
            I => \un114_pixel_6_1_5__un4_rowZ0Z_7_cascade_\
        );

    \I__1972\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10961\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__10961\,
            I => \N__10958\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__10958\,
            I => \un114_pixel_6_1_5__un4_rowZ0Z_1\
        );

    \I__1969\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10952\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__1967\ : Span4Mux_h
    port map (
            O => \N__10949\,
            I => \N__10943\
        );

    \I__1966\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10938\
        );

    \I__1965\ : InMux
    port map (
            O => \N__10947\,
            I => \N__10938\
        );

    \I__1964\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10935\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__10943\,
            I => \beamY_i_2\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__10938\,
            I => \beamY_i_2\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__10935\,
            I => \beamY_i_2\
        );

    \I__1960\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10925\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__1958\ : Span4Mux_v
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__10919\,
            I => \un114_pixel_6_1_5__chessboardpixel_un200_pixellto4Z0Z_1\
        );

    \I__1956\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10910\
        );

    \I__1955\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10910\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__10910\,
            I => \N__10907\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__10907\,
            I => \N__10904\
        );

    \I__1952\ : Span4Mux_h
    port map (
            O => \N__10904\,
            I => \N__10900\
        );

    \I__1951\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10897\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__10900\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__10897\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0\
        );

    \I__1948\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__1946\ : Span12Mux_s9_v
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__1945\ : Odrv12
    port map (
            O => \N__10883\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4OZ0\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__10880\,
            I => \chessboardpixel_un200_pixellt10_cascade_\
        );

    \I__1943\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10874\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__1941\ : Span4Mux_h
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__10868\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5
        );

    \I__1939\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__10862\,
            I => \N__10856\
        );

    \I__1937\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10846\
        );

    \I__1936\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10846\
        );

    \I__1935\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10846\
        );

    \I__1934\ : Span4Mux_h
    port map (
            O => \N__10856\,
            I => \N__10843\
        );

    \I__1933\ : InMux
    port map (
            O => \N__10855\,
            I => \N__10838\
        );

    \I__1932\ : InMux
    port map (
            O => \N__10854\,
            I => \N__10838\
        );

    \I__1931\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10835\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10832\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__10843\,
            I => chary_if_generate_plus_mult1_un68_sum_c5_0
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__10838\,
            I => chary_if_generate_plus_mult1_un68_sum_c5_0
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__10835\,
            I => chary_if_generate_plus_mult1_un68_sum_c5_0
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__10832\,
            I => chary_if_generate_plus_mult1_un68_sum_c5_0
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__10823\,
            I => \chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_cascade_\
        );

    \I__1924\ : InMux
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__10817\,
            I => \un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1Z0Z_1\
        );

    \I__1922\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__10811\,
            I => \N__10807\
        );

    \I__1920\ : InMux
    port map (
            O => \N__10810\,
            I => \N__10804\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__10807\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__10804\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__1916\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10793\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__10793\,
            I => \N__10790\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__10790\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0\
        );

    \I__1913\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10784\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__10784\,
            I => un4_beamy_0
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__10781\,
            I => \un13_beamylt10_0_cascade_\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1909\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10768\
        );

    \I__1908\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10765\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__10773\,
            I => \N__10762\
        );

    \I__1906\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10759\
        );

    \I__1905\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10756\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__10768\,
            I => \N__10751\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__10765\,
            I => \N__10751\
        );

    \I__1902\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10748\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__10759\,
            I => \beamXZ0Z_4\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__10756\,
            I => \beamXZ0Z_4\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__10751\,
            I => \beamXZ0Z_4\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__10748\,
            I => \beamXZ0Z_4\
        );

    \I__1897\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10732\
        );

    \I__1896\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10729\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__10737\,
            I => \N__10726\
        );

    \I__1894\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10723\
        );

    \I__1893\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10720\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__10732\,
            I => \N__10715\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__10729\,
            I => \N__10715\
        );

    \I__1890\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10712\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__10723\,
            I => \beamXZ0Z_3\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__10720\,
            I => \beamXZ0Z_3\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__10715\,
            I => \beamXZ0Z_3\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__10712\,
            I => \beamXZ0Z_3\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__1884\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__10697\,
            I => un18_beamylt5_0
        );

    \I__1882\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__10691\,
            I => \N__10683\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__10690\,
            I => \N__10680\
        );

    \I__1879\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10675\
        );

    \I__1878\ : InMux
    port map (
            O => \N__10688\,
            I => \N__10675\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__10687\,
            I => \N__10672\
        );

    \I__1876\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10669\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__10683\,
            I => \N__10666\
        );

    \I__1874\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10663\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__10675\,
            I => \N__10660\
        );

    \I__1872\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10657\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__10669\,
            I => \beamXZ0Z_5\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__10666\,
            I => \beamXZ0Z_5\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__10663\,
            I => \beamXZ0Z_5\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__10660\,
            I => \beamXZ0Z_5\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__10657\,
            I => \beamXZ0Z_5\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__10646\,
            I => \un18_beamylt5_0_cascade_\
        );

    \I__1865\ : InMux
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__10640\,
            I => \un114_pixel_6_1_5__un15_beamyZ0Z_0\
        );

    \I__1863\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10630\
        );

    \I__1862\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10627\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__10635\,
            I => \N__10624\
        );

    \I__1860\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10621\
        );

    \I__1859\ : InMux
    port map (
            O => \N__10633\,
            I => \N__10618\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__10630\,
            I => \N__10613\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__10627\,
            I => \N__10613\
        );

    \I__1856\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10610\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__10621\,
            I => \beamXZ0Z_8\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__10618\,
            I => \beamXZ0Z_8\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__10613\,
            I => \beamXZ0Z_8\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__10610\,
            I => \beamXZ0Z_8\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__10601\,
            I => \N__10595\
        );

    \I__1850\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10591\
        );

    \I__1849\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10588\
        );

    \I__1848\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10585\
        );

    \I__1847\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10582\
        );

    \I__1846\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10579\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__10591\,
            I => \beamXZ0Z_9\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__10588\,
            I => \beamXZ0Z_9\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__10585\,
            I => \beamXZ0Z_9\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__10582\,
            I => \beamXZ0Z_9\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__10579\,
            I => \beamXZ0Z_9\
        );

    \I__1840\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10560\
        );

    \I__1839\ : InMux
    port map (
            O => \N__10567\,
            I => \N__10555\
        );

    \I__1838\ : InMux
    port map (
            O => \N__10566\,
            I => \N__10555\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__10565\,
            I => \N__10552\
        );

    \I__1836\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10549\
        );

    \I__1835\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10546\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__10560\,
            I => \N__10541\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__10555\,
            I => \N__10541\
        );

    \I__1832\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10538\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__10549\,
            I => \beamXZ0Z_6\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__10546\,
            I => \beamXZ0Z_6\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__10541\,
            I => \beamXZ0Z_6\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__10538\,
            I => \beamXZ0Z_6\
        );

    \I__1827\ : InMux
    port map (
            O => \N__10529\,
            I => \N__10526\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__10526\,
            I => \un114_pixel_6_1_5__un18_beamylto9Z0Z_2\
        );

    \I__1825\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10520\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__10520\,
            I => \N__10514\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__10519\,
            I => \N__10511\
        );

    \I__1822\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10508\
        );

    \I__1821\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10505\
        );

    \I__1820\ : Span4Mux_v
    port map (
            O => \N__10514\,
            I => \N__10502\
        );

    \I__1819\ : InMux
    port map (
            O => \N__10511\,
            I => \N__10499\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__10508\,
            I => \beamXZ0Z_2\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__10505\,
            I => \beamXZ0Z_2\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__10502\,
            I => \beamXZ0Z_2\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__10499\,
            I => \beamXZ0Z_2\
        );

    \I__1814\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10483\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__10489\,
            I => \N__10480\
        );

    \I__1812\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10477\
        );

    \I__1811\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10474\
        );

    \I__1810\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10471\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__10483\,
            I => \N__10468\
        );

    \I__1808\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10465\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__10477\,
            I => \beamXZ0Z_1\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__10474\,
            I => \beamXZ0Z_1\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__10471\,
            I => \beamXZ0Z_1\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__10468\,
            I => \beamXZ0Z_1\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__10465\,
            I => \beamXZ0Z_1\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__1801\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__10448\,
            I => \un114_pixel_6_1_5__un13_beamylto2Z0Z_0\
        );

    \I__1799\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10439\
        );

    \I__1798\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10439\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__10439\,
            I => \un114_pixel_6_1_5__un15_beamyZ0Z_1\
        );

    \I__1796\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__10433\,
            I => un4_beamy_0_0
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__10421\,
            I => \un114_pixel_6_1_5__g3_0_0_0\
        );

    \I__1790\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__10415\,
            I => un13_beamylt10_0
        );

    \I__1788\ : InMux
    port map (
            O => \N__10412\,
            I => \bfn_6_6_0_\
        );

    \I__1787\ : InMux
    port map (
            O => \N__10409\,
            I => un5_visiblex_cry_8
        );

    \I__1786\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10403\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__10403\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0\
        );

    \I__1784\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__10397\,
            I => \N__10393\
        );

    \I__1782\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10390\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__10393\,
            I => \N__10387\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__10390\,
            I => \N__10384\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__10387\,
            I => if_generate_plus_mult1_un54_sum_axbxc5
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__10384\,
            I => if_generate_plus_mult1_un54_sum_axbxc5
        );

    \I__1777\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__10373\,
            I => \N__10369\
        );

    \I__1774\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10366\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__10369\,
            I => if_generate_plus_mult1_un61_sum_axbxc5
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__10366\,
            I => if_generate_plus_mult1_un61_sum_axbxc5
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__10361\,
            I => \un114_pixel_6_1_5__un3_beamxZ0Z_5_cascade_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__10355\,
            I => \un114_pixel_6_1_5__un3_beamxZ0Z_7\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__1767\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__10346\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i
        );

    \I__1765\ : InMux
    port map (
            O => \N__10343\,
            I => un5_visiblex_cry_0
        );

    \I__1764\ : InMux
    port map (
            O => \N__10340\,
            I => un5_visiblex_cry_1
        );

    \I__1763\ : InMux
    port map (
            O => \N__10337\,
            I => un5_visiblex_cry_2
        );

    \I__1762\ : InMux
    port map (
            O => \N__10334\,
            I => un5_visiblex_cry_3
        );

    \I__1761\ : InMux
    port map (
            O => \N__10331\,
            I => un5_visiblex_cry_4
        );

    \I__1760\ : InMux
    port map (
            O => \N__10328\,
            I => un5_visiblex_cry_5
        );

    \I__1759\ : InMux
    port map (
            O => \N__10325\,
            I => un5_visiblex_cry_6
        );

    \I__1758\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10317\
        );

    \I__1757\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10314\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__10320\,
            I => \N__10311\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__10317\,
            I => \N__10307\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__10314\,
            I => \N__10302\
        );

    \I__1753\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10296\
        );

    \I__1752\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10296\
        );

    \I__1751\ : Span4Mux_s3_h
    port map (
            O => \N__10307\,
            I => \N__10292\
        );

    \I__1750\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10287\
        );

    \I__1749\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10287\
        );

    \I__1748\ : Span4Mux_s3_h
    port map (
            O => \N__10302\,
            I => \N__10284\
        );

    \I__1747\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10281\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__10296\,
            I => \N__10278\
        );

    \I__1745\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10275\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__10292\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__10287\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__10284\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__10281\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__10278\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__10275\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__10262\,
            I => \N__10254\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__10261\,
            I => \N__10250\
        );

    \I__1736\ : InMux
    port map (
            O => \N__10260\,
            I => \N__10244\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10244\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__10258\,
            I => \N__10234\
        );

    \I__1733\ : InMux
    port map (
            O => \N__10257\,
            I => \N__10231\
        );

    \I__1732\ : InMux
    port map (
            O => \N__10254\,
            I => \N__10228\
        );

    \I__1731\ : InMux
    port map (
            O => \N__10253\,
            I => \N__10225\
        );

    \I__1730\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10222\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__10249\,
            I => \N__10219\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__10244\,
            I => \N__10216\
        );

    \I__1727\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10213\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10208\
        );

    \I__1725\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10205\
        );

    \I__1724\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10200\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10200\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__10238\,
            I => \N__10195\
        );

    \I__1721\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10192\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10189\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__10231\,
            I => \N__10186\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10183\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10180\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N__10177\
        );

    \I__1715\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10174\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__10216\,
            I => \N__10169\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__10213\,
            I => \N__10169\
        );

    \I__1712\ : InMux
    port map (
            O => \N__10212\,
            I => \N__10166\
        );

    \I__1711\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10163\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__10208\,
            I => \N__10160\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__10205\,
            I => \N__10155\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__10200\,
            I => \N__10155\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10152\
        );

    \I__1706\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10147\
        );

    \I__1705\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10147\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__10192\,
            I => \N__10142\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__10189\,
            I => \N__10142\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__10186\,
            I => \N__10137\
        );

    \I__1701\ : Span4Mux_v
    port map (
            O => \N__10183\,
            I => \N__10137\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__10180\,
            I => \N__10128\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__10177\,
            I => \N__10128\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__10174\,
            I => \N__10128\
        );

    \I__1697\ : Span4Mux_s1_h
    port map (
            O => \N__10169\,
            I => \N__10128\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__10166\,
            I => \N__10119\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10163\,
            I => \N__10119\
        );

    \I__1694\ : Sp12to4
    port map (
            O => \N__10160\,
            I => \N__10119\
        );

    \I__1693\ : Span12Mux_s4_h
    port map (
            O => \N__10155\,
            I => \N__10119\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__10152\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__10147\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__10142\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__10137\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__10128\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1687\ : Odrv12
    port map (
            O => \N__10119\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__10106\,
            I => \N__10101\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__10105\,
            I => \N__10098\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10104\,
            I => \N__10091\
        );

    \I__1683\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10087\
        );

    \I__1682\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10084\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__10097\,
            I => \N__10081\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__10096\,
            I => \N__10078\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__10095\,
            I => \N__10075\
        );

    \I__1678\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10072\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__10091\,
            I => \N__10069\
        );

    \I__1676\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10066\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__10087\,
            I => \N__10063\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__10084\,
            I => \N__10060\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10057\
        );

    \I__1672\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10054\
        );

    \I__1671\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10051\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10044\
        );

    \I__1669\ : Span4Mux_v
    port map (
            O => \N__10069\,
            I => \N__10044\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__10066\,
            I => \N__10044\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__10063\,
            I => \N__10037\
        );

    \I__1666\ : Span4Mux_h
    port map (
            O => \N__10060\,
            I => \N__10037\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__10057\,
            I => \N__10037\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__10054\,
            I => \N__10034\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10051\,
            I => \N__10029\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__10044\,
            I => \N__10029\
        );

    \I__1661\ : Odrv4
    port map (
            O => \N__10037\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1660\ : Odrv4
    port map (
            O => \N__10034\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__10029\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1658\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10011\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10011\
        );

    \I__1656\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10008\
        );

    \I__1655\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10005\
        );

    \I__1654\ : InMux
    port map (
            O => \N__10018\,
            I => \N__10000\
        );

    \I__1653\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10000\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10016\,
            I => \N__9997\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__10011\,
            I => \N__9994\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__9989\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__10005\,
            I => \N__9989\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__10000\,
            I => \N__9981\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__9997\,
            I => \N__9976\
        );

    \I__1646\ : Span4Mux_h
    port map (
            O => \N__9994\,
            I => \N__9976\
        );

    \I__1645\ : Span4Mux_h
    port map (
            O => \N__9989\,
            I => \N__9973\
        );

    \I__1644\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9962\
        );

    \I__1643\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9962\
        );

    \I__1642\ : InMux
    port map (
            O => \N__9986\,
            I => \N__9962\
        );

    \I__1641\ : InMux
    port map (
            O => \N__9985\,
            I => \N__9962\
        );

    \I__1640\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9962\
        );

    \I__1639\ : Odrv12
    port map (
            O => \N__9981\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__9976\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__9973\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__9962\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__1635\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9948\
        );

    \I__1634\ : InMux
    port map (
            O => \N__9952\,
            I => \N__9943\
        );

    \I__1633\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9943\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__9948\,
            I => chary_if_generate_plus_mult1_un68_sum_ac0_5
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__9943\,
            I => chary_if_generate_plus_mult1_un68_sum_ac0_5
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__9938\,
            I => \chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_\
        );

    \I__1629\ : InMux
    port map (
            O => \N__9935\,
            I => \N__9932\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__9932\,
            I => \beamY_RNIL0E2QG2Z0Z_3\
        );

    \I__1627\ : InMux
    port map (
            O => \N__9929\,
            I => \N__9926\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__9926\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93\
        );

    \I__1625\ : InMux
    port map (
            O => \N__9923\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__9920\,
            I => \N__9917\
        );

    \I__1623\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9914\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__9914\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4\
        );

    \I__1621\ : InMux
    port map (
            O => \N__9911\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__1620\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__9905\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__1618\ : InMux
    port map (
            O => \N__9902\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__1617\ : InMux
    port map (
            O => \N__9899\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__9896\,
            I => \N__9892\
        );

    \I__1615\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9888\
        );

    \I__1614\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9883\
        );

    \I__1613\ : InMux
    port map (
            O => \N__9891\,
            I => \N__9883\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__9888\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__9883\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__1609\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__9872\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i
        );

    \I__1607\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9863\
        );

    \I__1606\ : InMux
    port map (
            O => \N__9868\,
            I => \N__9863\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__9863\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__1604\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__9857\,
            I => g1
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__9854\,
            I => \N__9848\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__9853\,
            I => \N__9840\
        );

    \I__1600\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9836\
        );

    \I__1599\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9833\
        );

    \I__1598\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9830\
        );

    \I__1597\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9827\
        );

    \I__1596\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9822\
        );

    \I__1595\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9822\
        );

    \I__1594\ : InMux
    port map (
            O => \N__9844\,
            I => \N__9817\
        );

    \I__1593\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9817\
        );

    \I__1592\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9814\
        );

    \I__1591\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9811\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9808\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__9833\,
            I => \N__9799\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__9830\,
            I => \N__9799\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__9827\,
            I => \N__9799\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__9822\,
            I => \N__9799\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__9817\,
            I => \N__9793\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__9814\,
            I => \N__9793\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__9811\,
            I => \N__9790\
        );

    \I__1582\ : Span4Mux_v
    port map (
            O => \N__9808\,
            I => \N__9785\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__9799\,
            I => \N__9785\
        );

    \I__1580\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9782\
        );

    \I__1579\ : Span4Mux_h
    port map (
            O => \N__9793\,
            I => \N__9779\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__9790\,
            I => \beamYZ0Z_4\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__9785\,
            I => \beamYZ0Z_4\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__9782\,
            I => \beamYZ0Z_4\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__9779\,
            I => \beamYZ0Z_4\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__9770\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cascade_\
        );

    \I__1573\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9764\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__9764\,
            I => m511_0_x2_1_2
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__9761\,
            I => \G_7_0_m2_1_1_1_cascade_\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__9758\,
            I => \G_7_0_m2_1_1_cascade_\
        );

    \I__1569\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__9752\,
            I => \G_7_0_m2_1_0\
        );

    \I__1567\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9739\
        );

    \I__1566\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9739\
        );

    \I__1565\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9739\
        );

    \I__1564\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9736\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__9739\,
            I => \N__9733\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__9736\,
            I => \N__9730\
        );

    \I__1561\ : Span4Mux_h
    port map (
            O => \N__9733\,
            I => \N__9727\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__9730\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__9727\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__1558\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9718\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__9721\,
            I => \N__9714\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__9718\,
            I => \N__9710\
        );

    \I__1555\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9707\
        );

    \I__1554\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9702\
        );

    \I__1553\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9702\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__9710\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__9707\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__9702\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__9695\,
            I => \un114_pixel_6_1_5__g0_1Z0Z_4_cascade_\
        );

    \I__1548\ : InMux
    port map (
            O => \N__9692\,
            I => \N__9685\
        );

    \I__1547\ : InMux
    port map (
            O => \N__9691\,
            I => \N__9682\
        );

    \I__1546\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9677\
        );

    \I__1545\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9677\
        );

    \I__1544\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9674\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__9685\,
            I => \N__9665\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__9682\,
            I => \N__9665\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__9677\,
            I => \N__9660\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__9674\,
            I => \N__9660\
        );

    \I__1539\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9657\
        );

    \I__1538\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9654\
        );

    \I__1537\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9651\
        );

    \I__1536\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9648\
        );

    \I__1535\ : Span4Mux_v
    port map (
            O => \N__9665\,
            I => \N__9645\
        );

    \I__1534\ : Span4Mux_v
    port map (
            O => \N__9660\,
            I => \N__9640\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__9657\,
            I => \N__9640\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__9654\,
            I => \N__9637\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__9651\,
            I => \beamYZ0Z_5\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__9648\,
            I => \beamYZ0Z_5\
        );

    \I__1529\ : Odrv4
    port map (
            O => \N__9645\,
            I => \beamYZ0Z_5\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__9640\,
            I => \beamYZ0Z_5\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__9637\,
            I => \beamYZ0Z_5\
        );

    \I__1526\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9620\
        );

    \I__1525\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9617\
        );

    \I__1524\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9610\
        );

    \I__1523\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9610\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__9620\,
            I => \N__9600\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__9617\,
            I => \N__9600\
        );

    \I__1520\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9595\
        );

    \I__1519\ : InMux
    port map (
            O => \N__9615\,
            I => \N__9595\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__9610\,
            I => \N__9592\
        );

    \I__1517\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9589\
        );

    \I__1516\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9585\
        );

    \I__1515\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9580\
        );

    \I__1514\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9580\
        );

    \I__1513\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9577\
        );

    \I__1512\ : Span4Mux_v
    port map (
            O => \N__9600\,
            I => \N__9574\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__9595\,
            I => \N__9567\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__9592\,
            I => \N__9567\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__9589\,
            I => \N__9567\
        );

    \I__1508\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9564\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__9585\,
            I => \N__9561\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__9580\,
            I => \N__9558\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__9577\,
            I => \N__9553\
        );

    \I__1504\ : Span4Mux_v
    port map (
            O => \N__9574\,
            I => \N__9553\
        );

    \I__1503\ : Span4Mux_h
    port map (
            O => \N__9567\,
            I => \N__9550\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__9564\,
            I => \N__9547\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__9561\,
            I => \N__9544\
        );

    \I__1500\ : Span4Mux_s2_h
    port map (
            O => \N__9558\,
            I => \N__9541\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__9553\,
            I => \beamYZ0Z_9\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__9550\,
            I => \beamYZ0Z_9\
        );

    \I__1497\ : Odrv12
    port map (
            O => \N__9547\,
            I => \beamYZ0Z_9\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__9544\,
            I => \beamYZ0Z_9\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__9541\,
            I => \beamYZ0Z_9\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__9530\,
            I => \N__9527\
        );

    \I__1493\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9516\
        );

    \I__1492\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9516\
        );

    \I__1491\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9511\
        );

    \I__1490\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9511\
        );

    \I__1489\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9507\
        );

    \I__1488\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9502\
        );

    \I__1487\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9502\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__9516\,
            I => \N__9496\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__9511\,
            I => \N__9493\
        );

    \I__1484\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9488\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9483\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__9502\,
            I => \N__9483\
        );

    \I__1481\ : InMux
    port map (
            O => \N__9501\,
            I => \N__9478\
        );

    \I__1480\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9473\
        );

    \I__1479\ : InMux
    port map (
            O => \N__9499\,
            I => \N__9473\
        );

    \I__1478\ : Span4Mux_v
    port map (
            O => \N__9496\,
            I => \N__9468\
        );

    \I__1477\ : Span4Mux_v
    port map (
            O => \N__9493\,
            I => \N__9468\
        );

    \I__1476\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9463\
        );

    \I__1475\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9463\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__9488\,
            I => \N__9460\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__9483\,
            I => \N__9457\
        );

    \I__1472\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9452\
        );

    \I__1471\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9452\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__9478\,
            I => \N__9447\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__9473\,
            I => \N__9447\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__9468\,
            I => \N__9442\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__9463\,
            I => \N__9442\
        );

    \I__1466\ : Odrv12
    port map (
            O => \N__9460\,
            I => \beamYZ0Z_7\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__9457\,
            I => \beamYZ0Z_7\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__9452\,
            I => \beamYZ0Z_7\
        );

    \I__1463\ : Odrv12
    port map (
            O => \N__9447\,
            I => \beamYZ0Z_7\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__9442\,
            I => \beamYZ0Z_7\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__9431\,
            I => \N__9427\
        );

    \I__1460\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9420\
        );

    \I__1459\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9420\
        );

    \I__1458\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9417\
        );

    \I__1457\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9414\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__9420\,
            I => \N__9402\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9402\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__9414\,
            I => \N__9402\
        );

    \I__1453\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9399\
        );

    \I__1452\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9396\
        );

    \I__1451\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9393\
        );

    \I__1450\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9390\
        );

    \I__1449\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9387\
        );

    \I__1448\ : Span4Mux_v
    port map (
            O => \N__9402\,
            I => \N__9382\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__9399\,
            I => \N__9382\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__9396\,
            I => \N__9377\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__9393\,
            I => \N__9377\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__9390\,
            I => \beamYZ0Z_6\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__9387\,
            I => \beamYZ0Z_6\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__9382\,
            I => \beamYZ0Z_6\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__9377\,
            I => \beamYZ0Z_6\
        );

    \I__1440\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9365\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__9362\,
            I => \un114_pixel_6_1_5__g0_0Z0Z_4\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__9359\,
            I => \un114_pixel_6_1_5__g0_0Z0Z_3_cascade_\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__9356\,
            I => \un114_pixel_6_1_5__g2_0Z0Z_0_cascade_\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__9353\,
            I => \N__9341\
        );

    \I__1434\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9337\
        );

    \I__1433\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9332\
        );

    \I__1432\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9329\
        );

    \I__1431\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9325\
        );

    \I__1430\ : InMux
    port map (
            O => \N__9348\,
            I => \N__9320\
        );

    \I__1429\ : InMux
    port map (
            O => \N__9347\,
            I => \N__9320\
        );

    \I__1428\ : InMux
    port map (
            O => \N__9346\,
            I => \N__9315\
        );

    \I__1427\ : InMux
    port map (
            O => \N__9345\,
            I => \N__9315\
        );

    \I__1426\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9310\
        );

    \I__1425\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9310\
        );

    \I__1424\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9307\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__9337\,
            I => \N__9304\
        );

    \I__1422\ : InMux
    port map (
            O => \N__9336\,
            I => \N__9299\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9299\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9290\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9290\
        );

    \I__1418\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9287\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__9325\,
            I => \N__9280\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__9320\,
            I => \N__9280\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9280\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__9310\,
            I => \N__9277\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__9307\,
            I => \N__9274\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__9304\,
            I => \N__9269\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__9299\,
            I => \N__9269\
        );

    \I__1410\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9262\
        );

    \I__1409\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9262\
        );

    \I__1408\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9262\
        );

    \I__1407\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9257\
        );

    \I__1406\ : Span4Mux_v
    port map (
            O => \N__9290\,
            I => \N__9248\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__9287\,
            I => \N__9248\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__9280\,
            I => \N__9248\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__9277\,
            I => \N__9248\
        );

    \I__1402\ : Span4Mux_v
    port map (
            O => \N__9274\,
            I => \N__9241\
        );

    \I__1401\ : Span4Mux_h
    port map (
            O => \N__9269\,
            I => \N__9241\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__9262\,
            I => \N__9241\
        );

    \I__1399\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9238\
        );

    \I__1398\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9235\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__9257\,
            I => \beamYZ0Z_8\
        );

    \I__1396\ : Odrv4
    port map (
            O => \N__9248\,
            I => \beamYZ0Z_8\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__9241\,
            I => \beamYZ0Z_8\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__9238\,
            I => \beamYZ0Z_8\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9235\,
            I => \beamYZ0Z_8\
        );

    \I__1392\ : InMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__9218\,
            I => \un114_pixel_6_1_5__g0_0_1Z0Z_1\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__9215\,
            I => \un114_pixel_6_1_5__un1_beamylto9Z0Z_0_cascade_\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__9212\,
            I => \un114_pixel_6_1_5__un1_beamylto9_3_cascade_\
        );

    \I__1387\ : IoInMux
    port map (
            O => \N__9209\,
            I => \N__9206\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__1385\ : IoSpan4Mux
    port map (
            O => \N__9203\,
            I => \N__9199\
        );

    \I__1384\ : IoInMux
    port map (
            O => \N__9202\,
            I => \N__9196\
        );

    \I__1383\ : Span4Mux_s0_v
    port map (
            O => \N__9199\,
            I => \N__9193\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__9196\,
            I => \N__9190\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__9193\,
            I => \N__9187\
        );

    \I__1380\ : Span4Mux_s3_v
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__1379\ : Span4Mux_v
    port map (
            O => \N__9187\,
            I => \N__9179\
        );

    \I__1378\ : Span4Mux_v
    port map (
            O => \N__9184\,
            I => \N__9179\
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__9179\,
            I => \VSync_c\
        );

    \I__1376\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9171\
        );

    \I__1375\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9166\
        );

    \I__1374\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9166\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__9171\,
            I => un8_beamy_3
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__9166\,
            I => un8_beamy_3
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__9161\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cascade_\
        );

    \I__1370\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__9152\,
            I => \N__9145\
        );

    \I__1367\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9142\
        );

    \I__1366\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9139\
        );

    \I__1365\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9134\
        );

    \I__1364\ : InMux
    port map (
            O => \N__9148\,
            I => \N__9134\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__9145\,
            I => row_1_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__9142\,
            I => row_1_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__9139\,
            I => row_1_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__9134\,
            I => row_1_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \row_1_if_generate_plus_mult1_un82_sum_axbxc5_3Z0Z_1_cascade_\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__9122\,
            I => \N__9117\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__9121\,
            I => \N__9113\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9106\
        );

    \I__1355\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9101\
        );

    \I__1354\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9098\
        );

    \I__1353\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9092\
        );

    \I__1352\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9085\
        );

    \I__1351\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9085\
        );

    \I__1350\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9085\
        );

    \I__1349\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9082\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__9106\,
            I => \N__9079\
        );

    \I__1347\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9076\
        );

    \I__1346\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9069\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__9101\,
            I => \N__9066\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9063\
        );

    \I__1343\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9055\
        );

    \I__1342\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9055\
        );

    \I__1341\ : InMux
    port map (
            O => \N__9095\,
            I => \N__9055\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9052\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9049\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9044\
        );

    \I__1337\ : Span4Mux_s3_h
    port map (
            O => \N__9079\,
            I => \N__9044\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9041\
        );

    \I__1335\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9032\
        );

    \I__1334\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9032\
        );

    \I__1333\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9032\
        );

    \I__1332\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9032\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__9069\,
            I => \N__9029\
        );

    \I__1330\ : Span4Mux_s2_h
    port map (
            O => \N__9066\,
            I => \N__9026\
        );

    \I__1329\ : Span4Mux_s2_h
    port map (
            O => \N__9063\,
            I => \N__9023\
        );

    \I__1328\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9020\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__9055\,
            I => \N__9017\
        );

    \I__1326\ : Span4Mux_h
    port map (
            O => \N__9052\,
            I => \N__9012\
        );

    \I__1325\ : Span4Mux_s3_h
    port map (
            O => \N__9049\,
            I => \N__9012\
        );

    \I__1324\ : Span4Mux_v
    port map (
            O => \N__9044\,
            I => \N__9003\
        );

    \I__1323\ : Span4Mux_s3_h
    port map (
            O => \N__9041\,
            I => \N__9003\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__9032\,
            I => \N__9003\
        );

    \I__1321\ : Span4Mux_s3_h
    port map (
            O => \N__9029\,
            I => \N__9003\
        );

    \I__1320\ : Span4Mux_v
    port map (
            O => \N__9026\,
            I => \N__8998\
        );

    \I__1319\ : Span4Mux_v
    port map (
            O => \N__9023\,
            I => \N__8998\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__9020\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1317\ : Odrv12
    port map (
            O => \N__9017\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1316\ : Odrv4
    port map (
            O => \N__9012\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__9003\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__8998\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__8987\,
            I => \N__8983\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__8986\,
            I => \N__8980\
        );

    \I__1311\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8975\
        );

    \I__1310\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8975\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__8975\,
            I => un4_beamylt8_0
        );

    \I__1308\ : InMux
    port map (
            O => \N__8972\,
            I => un8_beamx_cry_6
        );

    \I__1307\ : InMux
    port map (
            O => \N__8969\,
            I => un8_beamx_cry_7
        );

    \I__1306\ : InMux
    port map (
            O => \N__8966\,
            I => \bfn_5_7_0_\
        );

    \I__1305\ : InMux
    port map (
            O => \N__8963\,
            I => un8_beamx_cry_9
        );

    \I__1304\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8957\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__8957\,
            I => row_1_if_generate_plus_mult1_un82_sum_axb4_i
        );

    \I__1302\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8951\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__8948\,
            I => \un114_pixel_6_1_5__un8_beamylto9Z0Z_0\
        );

    \I__1299\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__8942\,
            I => \N__8939\
        );

    \I__1297\ : Span4Mux_h
    port map (
            O => \N__8939\,
            I => \N__8936\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__8936\,
            I => un8_beamylt9_0
        );

    \I__1295\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8930\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__8930\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__1293\ : InMux
    port map (
            O => \N__8927\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__8924\,
            I => \N__8920\
        );

    \I__1291\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8915\
        );

    \I__1290\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8908\
        );

    \I__1289\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8908\
        );

    \I__1288\ : InMux
    port map (
            O => \N__8918\,
            I => \N__8908\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__8915\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__8908\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\
        );

    \I__1285\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__8900\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1282\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__8891\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i
        );

    \I__1280\ : InMux
    port map (
            O => \N__8888\,
            I => un8_beamx_cry_1
        );

    \I__1279\ : InMux
    port map (
            O => \N__8885\,
            I => un8_beamx_cry_2
        );

    \I__1278\ : InMux
    port map (
            O => \N__8882\,
            I => un8_beamx_cry_3
        );

    \I__1277\ : InMux
    port map (
            O => \N__8879\,
            I => un8_beamx_cry_4
        );

    \I__1276\ : InMux
    port map (
            O => \N__8876\,
            I => un8_beamx_cry_5
        );

    \I__1275\ : InMux
    port map (
            O => \N__8873\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1274\ : InMux
    port map (
            O => \N__8870\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__1273\ : InMux
    port map (
            O => \N__8867\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__1272\ : InMux
    port map (
            O => \N__8864\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__1271\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8855\
        );

    \I__1270\ : InMux
    port map (
            O => \N__8860\,
            I => \N__8855\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__8855\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__1268\ : InMux
    port map (
            O => \N__8852\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__1267\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__8846\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6\
        );

    \I__1265\ : InMux
    port map (
            O => \N__8843\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1263\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__8834\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9\
        );

    \I__1261\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__8828\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0\
        );

    \I__1259\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8822\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1257\ : Odrv12
    port map (
            O => \N__8819\,
            I => g2_1
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \chary_if_generate_plus_mult1_un68_sum_c5_0_cascade_\
        );

    \I__1255\ : CascadeMux
    port map (
            O => \N__8813\,
            I => \chary_if_generate_plus_mult1_un1_sum_axbxc3_1_1_cascade_\
        );

    \I__1254\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8801\
        );

    \I__1253\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8801\
        );

    \I__1252\ : InMux
    port map (
            O => \N__8808\,
            I => \N__8798\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__8807\,
            I => \N__8795\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8806\,
            I => \N__8792\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8787\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__8798\,
            I => \N__8787\
        );

    \I__1247\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8783\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__8792\,
            I => \N__8780\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__8787\,
            I => \N__8777\
        );

    \I__1244\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8774\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__8783\,
            I => chary_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__8780\,
            I => chary_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__8777\,
            I => chary_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__8774\,
            I => chary_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1239\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8759\
        );

    \I__1238\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8759\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__8759\,
            I => \N__8756\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__8756\,
            I => chary_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i
        );

    \I__1235\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8749\
        );

    \I__1234\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8746\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__8749\,
            I => \N__8741\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__8746\,
            I => \N__8741\
        );

    \I__1231\ : Span4Mux_h
    port map (
            O => \N__8741\,
            I => \N__8737\
        );

    \I__1230\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8734\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__8737\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_0
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__8734\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_0
        );

    \I__1227\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__1225\ : Span4Mux_s3_h
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__8720\,
            I => chary_if_generate_plus_mult1_un68_sum_c5_0_0
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__8717\,
            I => \un114_pixel_6_1_5__g0_17Z0Z_1_cascade_\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__8711\,
            I => chary_if_generate_plus_mult1_un75_sum_0_5
        );

    \I__1220\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8705\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__8702\,
            I => chary_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__1216\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8692\
        );

    \I__1215\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8689\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__8692\,
            I => \N__8686\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__8689\,
            I => chary_if_generate_plus_mult1_un61_sum_c4
        );

    \I__1212\ : Odrv12
    port map (
            O => \N__8686\,
            I => chary_if_generate_plus_mult1_un61_sum_c4
        );

    \I__1211\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__8678\,
            I => g1_0_3
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__8675\,
            I => \N__8670\
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__8674\,
            I => \N__8667\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__8673\,
            I => \N__8664\
        );

    \I__1206\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8659\
        );

    \I__1205\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8659\
        );

    \I__1204\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8656\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__8659\,
            I => \N__8653\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__8656\,
            I => \N__8648\
        );

    \I__1201\ : Span4Mux_h
    port map (
            O => \N__8653\,
            I => \N__8645\
        );

    \I__1200\ : InMux
    port map (
            O => \N__8652\,
            I => \N__8640\
        );

    \I__1199\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8640\
        );

    \I__1198\ : Span4Mux_h
    port map (
            O => \N__8648\,
            I => \N__8637\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__8645\,
            I => un5_visibley_c5
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__8640\,
            I => un5_visibley_c5
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__8637\,
            I => un5_visibley_c5
        );

    \I__1194\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8627\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__8627\,
            I => \beamY_RNIP8FF1_2Z0Z_7\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__8624\,
            I => \un4_beamylt6_cascade_\
        );

    \I__1191\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8615\
        );

    \I__1190\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8615\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8610\
        );

    \I__1188\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8606\
        );

    \I__1187\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8603\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__8610\,
            I => \N__8600\
        );

    \I__1185\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8597\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__8606\,
            I => \N__8592\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__8603\,
            I => \N__8592\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__8600\,
            I => \N__8589\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__8597\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__8592\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__8589\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__1178\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8572\
        );

    \I__1177\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8572\
        );

    \I__1176\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8566\
        );

    \I__1175\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8566\
        );

    \I__1174\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8561\
        );

    \I__1173\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8561\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__8572\,
            I => \N__8558\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__8571\,
            I => \N__8553\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__8566\,
            I => \N__8547\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__8561\,
            I => \N__8547\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__8558\,
            I => \N__8544\
        );

    \I__1167\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8535\
        );

    \I__1166\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8535\
        );

    \I__1165\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8535\
        );

    \I__1164\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8535\
        );

    \I__1163\ : Odrv4
    port map (
            O => \N__8547\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1162\ : Odrv4
    port map (
            O => \N__8544\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__8535\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__8528\,
            I => \beamY_RNIB6AOI5_0Z0Z_5_cascade_\
        );

    \I__1159\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8518\
        );

    \I__1158\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8509\
        );

    \I__1157\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8509\
        );

    \I__1156\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8509\
        );

    \I__1155\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8509\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8506\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__8509\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_d
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__8506\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_d
        );

    \I__1151\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__1149\ : Span4Mux_v
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__8492\,
            I => un5_visibley_c2
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__8489\,
            I => \N__8483\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__8488\,
            I => \N__8476\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__8487\,
            I => \N__8472\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__8486\,
            I => \N__8468\
        );

    \I__1143\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8465\
        );

    \I__1142\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8458\
        );

    \I__1141\ : InMux
    port map (
            O => \N__8481\,
            I => \N__8455\
        );

    \I__1140\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8448\
        );

    \I__1139\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8448\
        );

    \I__1138\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8448\
        );

    \I__1137\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8443\
        );

    \I__1136\ : InMux
    port map (
            O => \N__8472\,
            I => \N__8443\
        );

    \I__1135\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8440\
        );

    \I__1134\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8437\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__8465\,
            I => \N__8434\
        );

    \I__1132\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8429\
        );

    \I__1131\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8429\
        );

    \I__1130\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8426\
        );

    \I__1129\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8423\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8420\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__8455\,
            I => \N__8417\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__8448\,
            I => \N__8414\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__8443\,
            I => \N__8411\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__8440\,
            I => \N__8404\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__8437\,
            I => \N__8404\
        );

    \I__1122\ : Span4Mux_s3_h
    port map (
            O => \N__8434\,
            I => \N__8404\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__8429\,
            I => \N__8401\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__8426\,
            I => \N__8398\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__8423\,
            I => \N__8395\
        );

    \I__1118\ : Span4Mux_s3_h
    port map (
            O => \N__8420\,
            I => \N__8392\
        );

    \I__1117\ : Span4Mux_s3_h
    port map (
            O => \N__8417\,
            I => \N__8389\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__8414\,
            I => \N__8386\
        );

    \I__1115\ : Span12Mux_s3_h
    port map (
            O => \N__8411\,
            I => \N__8383\
        );

    \I__1114\ : Span4Mux_v
    port map (
            O => \N__8404\,
            I => \N__8378\
        );

    \I__1113\ : Span4Mux_s3_h
    port map (
            O => \N__8401\,
            I => \N__8378\
        );

    \I__1112\ : Span12Mux_s10_v
    port map (
            O => \N__8398\,
            I => \N__8375\
        );

    \I__1111\ : Span4Mux_s3_h
    port map (
            O => \N__8395\,
            I => \N__8370\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__8392\,
            I => \N__8370\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__8389\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__8386\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1107\ : Odrv12
    port map (
            O => \N__8383\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__8378\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__8375\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__8370\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1103\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8351\
        );

    \I__1102\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8351\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__8351\,
            I => row_1_if_generate_plus_mult1_un75_sum_c5
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__8348\,
            I => \if_generate_plus_mult1_un82_sum_axb4_x1_cascade_\
        );

    \I__1099\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8342\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__8342\,
            I => if_generate_plus_mult1_un82_sum_axb4_x0
        );

    \I__1097\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__1095\ : Span4Mux_s1_h
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__8330\,
            I => \beamY_RNIP8FF1_0Z0Z_7\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__8327\,
            I => \un114_pixel_6_1_5__un5_beamxZ0Z_3_cascade_\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__8324\,
            I => \un114_pixel_6_1_5__un5_beamxZ0Z_5_cascade_\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__8321\,
            I => \beamY_RNIP8FF1Z0Z_7_cascade_\
        );

    \I__1090\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8312\
        );

    \I__1089\ : InMux
    port map (
            O => \N__8317\,
            I => \N__8308\
        );

    \I__1088\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8303\
        );

    \I__1087\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8300\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__8312\,
            I => \N__8297\
        );

    \I__1085\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8294\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8291\
        );

    \I__1083\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8286\
        );

    \I__1082\ : InMux
    port map (
            O => \N__8306\,
            I => \N__8286\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__8303\,
            I => \N__8279\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8279\
        );

    \I__1079\ : Span4Mux_h
    port map (
            O => \N__8297\,
            I => \N__8279\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__8294\,
            I => un5_visibley_c6
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__8291\,
            I => un5_visibley_c6
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__8286\,
            I => un5_visibley_c6
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__8279\,
            I => un5_visibley_c6
        );

    \I__1074\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8264\
        );

    \I__1073\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8264\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__8264\,
            I => \N__8260\
        );

    \I__1071\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8257\
        );

    \I__1070\ : IoSpan4Mux
    port map (
            O => \N__8260\,
            I => \N__8252\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__8257\,
            I => \N__8252\
        );

    \I__1068\ : Span4Mux_s3_h
    port map (
            O => \N__8252\,
            I => \N__8249\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__8249\,
            I => chary_if_generate_plus_mult1_un40_sum_c4
        );

    \I__1066\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8243\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__8243\,
            I => \row_1_if_generate_plus_mult1_un61_sum_ac0_7_0Z0Z_1\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__8240\,
            I => \row_1_if_i4_mux_i_cascade_\
        );

    \I__1063\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8230\
        );

    \I__1062\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8225\
        );

    \I__1061\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8225\
        );

    \I__1060\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8220\
        );

    \I__1059\ : InMux
    port map (
            O => \N__8233\,
            I => \N__8220\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8230\,
            I => \N__8215\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__8225\,
            I => \N__8215\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__8220\,
            I => \N__8212\
        );

    \I__1055\ : Span4Mux_v
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__8212\,
            I => \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__8209\,
            I => \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\
        );

    \I__1052\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8201\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__8201\,
            I => row_1_if_i4_mux_i
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__8198\,
            I => \row_1_if_generate_plus_mult1_un75_sum_ac0_7_0Z0Z_1_cascade_\
        );

    \I__1049\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__8192\,
            I => \row_1_if_N_6\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__8189\,
            I => \if_generate_plus_mult1_un75_sum_axbxc3_cascade_\
        );

    \I__1046\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8182\
        );

    \I__1045\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8179\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__8182\,
            I => \N__8176\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__8179\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__8176\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__8171\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8165\,
            I => \N__8160\
        );

    \I__1038\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8155\
        );

    \I__1037\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8155\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__8160\,
            I => \N__8150\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__8155\,
            I => \N__8150\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__8150\,
            I => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0\
        );

    \I__1033\ : InMux
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8144\,
            I => if_generate_plus_mult1_un75_sum_axbxc3
        );

    \I__1031\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8138\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__8138\,
            I => \N__8134\
        );

    \I__1029\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1028\ : Span4Mux_v
    port map (
            O => \N__8134\,
            I => \N__8128\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__8128\,
            I => \un21_beamy_cry_7_c_RNIM7EZ0Z3\
        );

    \I__1025\ : Odrv12
    port map (
            O => \N__8125\,
            I => \un21_beamy_cry_7_c_RNIM7EZ0Z3\
        );

    \I__1024\ : InMux
    port map (
            O => \N__8120\,
            I => un21_beamy_cry_7
        );

    \I__1023\ : InMux
    port map (
            O => \N__8117\,
            I => \bfn_2_13_0_\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \if_generate_plus_mult1_un61_sum_axbxc5_cascade_\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__8111\,
            I => \N__8107\
        );

    \I__1020\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8104\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8101\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8104\,
            I => \row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__8101\,
            I => \row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__8096\,
            I => \row_1_if_generate_plus_mult1_un61_sum_ac0_7_dZ0_cascade_\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__8093\,
            I => \row_1_if_generate_plus_mult1_un61_sum_c5_cascade_\
        );

    \I__1014\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8084\
        );

    \I__1013\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8084\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1011\ : Odrv12
    port map (
            O => \N__8081\,
            I => row_1_if_generate_plus_mult1_un61_sum_axb4_i
        );

    \I__1010\ : CascadeMux
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1009\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8072\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8069\
        );

    \I__1007\ : Odrv12
    port map (
            O => \N__8069\,
            I => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_6\
        );

    \I__1006\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8060\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8060\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8060\,
            I => \N__8057\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__8057\,
            I => \un21_beamy_cry_1_c_RNIALZ0Z73\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8054\,
            I => un21_beamy_cry_1
        );

    \I__1001\ : InMux
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__8048\,
            I => \N__8044\
        );

    \I__999\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8041\
        );

    \I__998\ : Span4Mux_v
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__8038\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__995\ : Odrv12
    port map (
            O => \N__8035\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__994\ : InMux
    port map (
            O => \N__8030\,
            I => un21_beamy_cry_2
        );

    \I__993\ : InMux
    port map (
            O => \N__8027\,
            I => \N__8023\
        );

    \I__992\ : InMux
    port map (
            O => \N__8026\,
            I => \N__8020\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__8023\,
            I => \N__8017\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__8020\,
            I => \N__8014\
        );

    \I__989\ : Odrv12
    port map (
            O => \N__8017\,
            I => \un21_beamy_cry_3_c_RNIERZ0Z93\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__8014\,
            I => \un21_beamy_cry_3_c_RNIERZ0Z93\
        );

    \I__987\ : InMux
    port map (
            O => \N__8009\,
            I => un21_beamy_cry_3
        );

    \I__986\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8003\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__8003\,
            I => \N__7999\
        );

    \I__984\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__983\ : Odrv12
    port map (
            O => \N__7999\,
            I => \un21_beamy_cry_4_c_RNIGUAZ0Z3\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__7996\,
            I => \un21_beamy_cry_4_c_RNIGUAZ0Z3\
        );

    \I__981\ : InMux
    port map (
            O => \N__7991\,
            I => un21_beamy_cry_4
        );

    \I__980\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7985\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7981\
        );

    \I__978\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7978\
        );

    \I__977\ : Odrv12
    port map (
            O => \N__7981\,
            I => \un21_beamy_cry_5_c_RNII1CZ0Z3\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__7978\,
            I => \un21_beamy_cry_5_c_RNII1CZ0Z3\
        );

    \I__975\ : InMux
    port map (
            O => \N__7973\,
            I => un21_beamy_cry_5
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__973\ : InMux
    port map (
            O => \N__7967\,
            I => \N__7961\
        );

    \I__972\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7961\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__970\ : Odrv12
    port map (
            O => \N__7958\,
            I => \un21_beamy_cry_6_c_RNIK4DZ0Z3\
        );

    \I__969\ : InMux
    port map (
            O => \N__7955\,
            I => un21_beamy_cry_6
        );

    \I__968\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7948\
        );

    \I__967\ : InMux
    port map (
            O => \N__7951\,
            I => \N__7945\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__7948\,
            I => \beamY_fastZ0Z_7\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__7945\,
            I => \beamY_fastZ0Z_7\
        );

    \I__964\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7932\
        );

    \I__963\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7932\
        );

    \I__962\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7929\
        );

    \I__961\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7926\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__7932\,
            I => \beamY_fastZ0Z_6\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__7929\,
            I => \beamY_fastZ0Z_6\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__7926\,
            I => \beamY_fastZ0Z_6\
        );

    \I__957\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7910\
        );

    \I__956\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7910\
        );

    \I__955\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7910\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__7910\,
            I => \beamY_fastZ0Z_5\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__7907\,
            I => \un5_visibley_ac0_11_0_1_cascade_\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__7904\,
            I => \N__7900\
        );

    \I__951\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7896\
        );

    \I__950\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7891\
        );

    \I__949\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7891\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__7896\,
            I => \beamY_fastZ0Z_4\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__7891\,
            I => \beamY_fastZ0Z_4\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__7886\,
            I => \N__7882\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__7885\,
            I => \N__7879\
        );

    \I__944\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7874\
        );

    \I__943\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7874\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__7874\,
            I => \beamY_fastZ0Z_8\
        );

    \I__941\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__7868\,
            I => un5_visibley_c7
        );

    \I__939\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7862\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7856\
        );

    \I__937\ : InMux
    port map (
            O => \N__7861\,
            I => \N__7853\
        );

    \I__936\ : InMux
    port map (
            O => \N__7860\,
            I => \N__7850\
        );

    \I__935\ : InMux
    port map (
            O => \N__7859\,
            I => \N__7847\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__7856\,
            I => \beamY_fastZ0Z_3\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7853\,
            I => \beamY_fastZ0Z_3\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__7850\,
            I => \beamY_fastZ0Z_3\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__7847\,
            I => \beamY_fastZ0Z_3\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__7838\,
            I => \un5_visibley_c2_cascade_\
        );

    \I__929\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7829\
        );

    \I__928\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7826\
        );

    \I__927\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7821\
        );

    \I__926\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7821\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__7829\,
            I => \beamY_fastZ0Z_2\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__7826\,
            I => \beamY_fastZ0Z_2\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__7821\,
            I => \beamY_fastZ0Z_2\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__7814\,
            I => \beamY_fast_RNIT5UFZ0Z_4_cascade_\
        );

    \I__921\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__7808\,
            I => un5_visibley_ac0_7
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__7805\,
            I => \un5_visibley_ac0_7_cascade_\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__917\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7796\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__7796\,
            I => \N__7792\
        );

    \I__915\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7789\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__7792\,
            I => chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux
        );

    \I__913\ : LocalMux
    port map (
            O => \N__7789\,
            I => chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux
        );

    \I__912\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7781\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__7781\,
            I => \N__7778\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__7778\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__909\ : CascadeMux
    port map (
            O => \N__7775\,
            I => \N__7772\
        );

    \I__908\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7766\
        );

    \I__907\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7766\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__7766\,
            I => \N__7763\
        );

    \I__905\ : Span4Mux_v
    port map (
            O => \N__7763\,
            I => \N__7760\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__7760\,
            I => chary_if_generate_plus_mult1_un47_sum_axb3
        );

    \I__903\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7751\
        );

    \I__902\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7751\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__7751\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NEZ0\
        );

    \I__900\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7742\
        );

    \I__899\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7742\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__7742\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATKZ0\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__7739\,
            I => \beamY_i_2_cascade_\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__7736\,
            I => \N__7733\
        );

    \I__895\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7730\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__7730\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6UZ0\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__7727\,
            I => \N__7724\
        );

    \I__892\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__7721\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVHZ0Z1\
        );

    \I__890\ : InMux
    port map (
            O => \N__7718\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__889\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__7712\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEAZ0Z1\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__7709\,
            I => \N__7706\
        );

    \I__886\ : InMux
    port map (
            O => \N__7706\,
            I => \N__7703\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__7703\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8UZ0Z1\
        );

    \I__884\ : InMux
    port map (
            O => \N__7700\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__7697\,
            I => \N__7694\
        );

    \I__882\ : InMux
    port map (
            O => \N__7694\,
            I => \N__7691\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__7691\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HAZ0Z1\
        );

    \I__880\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__7685\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__878\ : InMux
    port map (
            O => \N__7682\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__877\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7674\
        );

    \I__876\ : InMux
    port map (
            O => \N__7678\,
            I => \N__7669\
        );

    \I__875\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7669\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__7674\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__873\ : LocalMux
    port map (
            O => \N__7669\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__871\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__7658\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__869\ : InMux
    port map (
            O => \N__7655\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__7652\,
            I => \N__7647\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__7651\,
            I => \N__7643\
        );

    \I__866\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7631\
        );

    \I__865\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7631\
        );

    \I__864\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7631\
        );

    \I__863\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7631\
        );

    \I__862\ : InMux
    port map (
            O => \N__7642\,
            I => \N__7631\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__7631\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9\
        );

    \I__860\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7625\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__7625\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__7622\,
            I => \N__7618\
        );

    \I__857\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7608\
        );

    \I__856\ : InMux
    port map (
            O => \N__7618\,
            I => \N__7608\
        );

    \I__855\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7608\
        );

    \I__854\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7603\
        );

    \I__853\ : InMux
    port map (
            O => \N__7615\,
            I => \N__7603\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7608\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__7603\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\
        );

    \I__850\ : InMux
    port map (
            O => \N__7598\,
            I => \N__7595\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__7595\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7
        );

    \I__848\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__7586\,
            I => if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx
        );

    \I__845\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7580\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__7580\,
            I => \beamY_RNIUUEM_0Z0Z_8\
        );

    \I__843\ : InMux
    port map (
            O => \N__7577\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__842\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__7571\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVLZ0Z21\
        );

    \I__840\ : InMux
    port map (
            O => \N__7568\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__839\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7562\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__7562\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1NZ0Z21\
        );

    \I__837\ : InMux
    port map (
            O => \N__7559\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__836\ : InMux
    port map (
            O => \N__7556\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__835\ : InMux
    port map (
            O => \N__7553\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__834\ : InMux
    port map (
            O => \N__7550\,
            I => \N__7544\
        );

    \I__833\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7544\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__7544\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__831\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__7538\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0\
        );

    \I__829\ : InMux
    port map (
            O => \N__7535\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__7532\,
            I => \chary_if_generate_plus_mult1_un61_sum_axb4_i_cascade_\
        );

    \I__827\ : InMux
    port map (
            O => \N__7529\,
            I => \N__7526\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__7526\,
            I => \un114_pixel_6_1_5__g0Z0Z_2\
        );

    \I__825\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7517\
        );

    \I__824\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7517\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__822\ : Odrv4
    port map (
            O => \N__7514\,
            I => chary_if_generate_plus_mult1_un61_sum_axb4_0
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__7511\,
            I => \chary_if_generate_plus_mult1_un61_sum_c4_cascade_\
        );

    \I__820\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7505\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__7505\,
            I => \N__7500\
        );

    \I__818\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7497\
        );

    \I__817\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7494\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__7500\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0
        );

    \I__815\ : LocalMux
    port map (
            O => \N__7497\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0
        );

    \I__814\ : LocalMux
    port map (
            O => \N__7494\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__7487\,
            I => \beamY_RNISDTA58Z0Z_5_cascade_\
        );

    \I__812\ : InMux
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__7481\,
            I => \beamY_RNIJ0797KZ0Z_4\
        );

    \I__810\ : InMux
    port map (
            O => \N__7478\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__809\ : InMux
    port map (
            O => \N__7475\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__808\ : InMux
    port map (
            O => \N__7472\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__807\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__7466\,
            I => \beamY_RNI2B511_0Z0Z_9\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__804\ : InMux
    port map (
            O => \N__7460\,
            I => \N__7457\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__7457\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_0
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__7454\,
            I => \chary_if_generate_plus_mult1_un68_sum_axb4_0_cascade_\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__7451\,
            I => \chary_if_generate_plus_mult1_un68_sum_axb4_i_cascade_\
        );

    \I__800\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__7445\,
            I => g1_0_2
        );

    \I__798\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7436\
        );

    \I__797\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7436\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__7436\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__794\ : InMux
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__7427\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_0
        );

    \I__792\ : InMux
    port map (
            O => \N__7424\,
            I => \N__7421\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__7421\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4_i_0
        );

    \I__790\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__7415\,
            I => g1_1
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__7412\,
            I => \g2_0_cascade_\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__7409\,
            I => \beamY_RNIV5SUC3_0Z0Z_9_cascade_\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__7406\,
            I => \N__7403\
        );

    \I__785\ : InMux
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__7400\,
            I => chary_if_generate_plus_mult1_un61_sum_axb4_0_1
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__7397\,
            I => \chary_if_generate_plus_mult1_un61_sum_axb4_0_cascade_\
        );

    \I__782\ : InMux
    port map (
            O => \N__7394\,
            I => \N__7385\
        );

    \I__781\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7385\
        );

    \I__780\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7382\
        );

    \I__779\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7377\
        );

    \I__778\ : InMux
    port map (
            O => \N__7390\,
            I => \N__7377\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__7385\,
            I => \beamY_RNIVADQVZ0Z_8\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__7382\,
            I => \beamY_RNIVADQVZ0Z_8\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__7377\,
            I => \beamY_RNIVADQVZ0Z_8\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__7370\,
            I => \N__7364\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__7369\,
            I => \N__7361\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__7368\,
            I => \N__7357\
        );

    \I__771\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7350\
        );

    \I__770\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7350\
        );

    \I__769\ : InMux
    port map (
            O => \N__7361\,
            I => \N__7350\
        );

    \I__768\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7345\
        );

    \I__767\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7345\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__7350\,
            I => \N__7342\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__7345\,
            I => \N__7339\
        );

    \I__764\ : Odrv12
    port map (
            O => \N__7342\,
            I => chary_if_generate_plus_mult1_un47_sum_c4
        );

    \I__763\ : Odrv4
    port map (
            O => \N__7339\,
            I => chary_if_generate_plus_mult1_un47_sum_c4
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__7334\,
            I => \N__7327\
        );

    \I__761\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7319\
        );

    \I__760\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7319\
        );

    \I__759\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7319\
        );

    \I__758\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7312\
        );

    \I__757\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7312\
        );

    \I__756\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7312\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__7319\,
            I => \N__7308\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__7312\,
            I => \N__7305\
        );

    \I__753\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7302\
        );

    \I__752\ : Odrv12
    port map (
            O => \N__7308\,
            I => chary_if_generate_plus_mult1_un47_sum_axb4
        );

    \I__751\ : Odrv4
    port map (
            O => \N__7305\,
            I => chary_if_generate_plus_mult1_un47_sum_axb4
        );

    \I__750\ : LocalMux
    port map (
            O => \N__7302\,
            I => chary_if_generate_plus_mult1_un47_sum_axb4
        );

    \I__749\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7292\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__7292\,
            I => \beamY_RNIV5SUC3Z0Z_9\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__7289\,
            I => \chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_cascade_\
        );

    \I__746\ : InMux
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__7283\,
            I => \beamY_RNIP8FF1_1Z0Z_7\
        );

    \I__744\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7275\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__7279\,
            I => \N__7271\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__7278\,
            I => \N__7265\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__7275\,
            I => \N__7262\
        );

    \I__740\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7257\
        );

    \I__739\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7257\
        );

    \I__738\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7254\
        );

    \I__737\ : InMux
    port map (
            O => \N__7269\,
            I => \N__7249\
        );

    \I__736\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7249\
        );

    \I__735\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7246\
        );

    \I__734\ : Odrv4
    port map (
            O => \N__7262\,
            I => \beamY_RNI93821Z0Z_9\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__7257\,
            I => \beamY_RNI93821Z0Z_9\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__7254\,
            I => \beamY_RNI93821Z0Z_9\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__7249\,
            I => \beamY_RNI93821Z0Z_9\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__7246\,
            I => \beamY_RNI93821Z0Z_9\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__7235\,
            I => \beamY_RNIBV5E51Z0Z_8_cascade_\
        );

    \I__728\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__7229\,
            I => \beamY_RNIBV5E51_0Z0Z_8\
        );

    \I__726\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7216\
        );

    \I__725\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7216\
        );

    \I__724\ : InMux
    port map (
            O => \N__7224\,
            I => \N__7216\
        );

    \I__723\ : InMux
    port map (
            O => \N__7223\,
            I => \N__7213\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__7216\,
            I => \N__7208\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__7213\,
            I => \N__7208\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__7208\,
            I => chary_if_generate_plus_mult1_un47_sum_axbxc5_2
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__7205\,
            I => \N__7200\
        );

    \I__718\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7190\
        );

    \I__717\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7190\
        );

    \I__716\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7190\
        );

    \I__715\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7190\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__7190\,
            I => \N__7186\
        );

    \I__713\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7183\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__7186\,
            I => chary_if_generate_plus_mult1_un47_sum_c5
        );

    \I__711\ : LocalMux
    port map (
            O => \N__7183\,
            I => chary_if_generate_plus_mult1_un47_sum_c5
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__7178\,
            I => \beamY_RNIVADQVZ0Z_8_cascade_\
        );

    \I__709\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7169\
        );

    \I__708\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7169\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__7169\,
            I => chary_if_generate_plus_mult1_un54_sum_ac0_5
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__7166\,
            I => \beamY_RNI93821Z0Z_9_cascade_\
        );

    \I__705\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7160\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__7160\,
            I => \beamY_RNIM5433_0Z0Z_8\
        );

    \I__703\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__7154\,
            I => \beamY_RNIIR4K3_0Z0Z_7\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__7151\,
            I => \beamY_RNIIR4K3_0Z0Z_7_cascade_\
        );

    \I__700\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7145\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__7145\,
            I => \beamY_RNIKM9GC_0Z0Z_9\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__7142\,
            I => \chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_\
        );

    \I__697\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7136\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__695\ : Odrv12
    port map (
            O => \N__7133\,
            I => \beamY_RNI9DSP2_0Z0Z_8\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__7130\,
            I => \beamY_RNI41384Z0Z_7_cascade_\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__7127\,
            I => \chary_if_generate_plus_mult1_un54_sum_ac0_5_1_cascade_\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__7124\,
            I => \un8_beamylt9_0_cascade_\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__7121\,
            I => \N__7118\
        );

    \I__690\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7115\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__7115\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74AZ0\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__7112\,
            I => \N__7107\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__7111\,
            I => \N__7103\
        );

    \I__686\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7099\
        );

    \I__685\ : InMux
    port map (
            O => \N__7107\,
            I => \N__7090\
        );

    \I__684\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7090\
        );

    \I__683\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7090\
        );

    \I__682\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7090\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7099\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__7090\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0\
        );

    \I__679\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__7082\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7
        );

    \I__677\ : InMux
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__7076\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__675\ : InMux
    port map (
            O => \N__7073\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__674\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__7067\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__7064\,
            I => \chary_if_generate_plus_mult1_un47_sum_axb4_cascade_\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__7061\,
            I => \beamY_RNIKM9GCZ0Z_9_cascade_\
        );

    \I__670\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7055\,
            I => \beamY_RNIM5433Z0Z_8\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__667\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7046\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__7046\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PUZ0Z3\
        );

    \I__665\ : InMux
    port map (
            O => \N__7043\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__7040\,
            I => \N__7037\
        );

    \I__663\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__7034\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJZ0Z4\
        );

    \I__661\ : InMux
    port map (
            O => \N__7031\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__660\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__7025\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__658\ : InMux
    port map (
            O => \N__7022\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__7019\,
            I => \N__7014\
        );

    \I__656\ : InMux
    port map (
            O => \N__7018\,
            I => \N__7009\
        );

    \I__655\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7000\
        );

    \I__654\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7000\
        );

    \I__653\ : InMux
    port map (
            O => \N__7013\,
            I => \N__7000\
        );

    \I__652\ : InMux
    port map (
            O => \N__7012\,
            I => \N__7000\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__7009\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__7000\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5\
        );

    \I__649\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__6992\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__647\ : InMux
    port map (
            O => \N__6989\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__6986\,
            I => \N__6983\
        );

    \I__645\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6980\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__6977\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8AZ0Z6\
        );

    \I__642\ : InMux
    port map (
            O => \N__6974\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__641\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6968\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__6968\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RHZ0Z9\
        );

    \I__639\ : InMux
    port map (
            O => \N__6965\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__6962\,
            I => \N__6958\
        );

    \I__637\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6949\
        );

    \I__636\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6949\
        );

    \I__635\ : InMux
    port map (
            O => \N__6957\,
            I => \N__6949\
        );

    \I__634\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6946\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__6949\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__6946\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__6941\,
            I => \N__6938\
        );

    \I__630\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6935\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__6935\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1\
        );

    \I__628\ : InMux
    port map (
            O => \N__6932\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__627\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6926\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__6926\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRUZ0Z85\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__6923\,
            I => \N__6919\
        );

    \I__624\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6916\
        );

    \I__623\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6913\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__6916\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__6913\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2\
        );

    \I__620\ : InMux
    port map (
            O => \N__6908\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__619\ : InMux
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__6902\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__617\ : InMux
    port map (
            O => \N__6899\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__6896\,
            I => \N__6893\
        );

    \I__615\ : InMux
    port map (
            O => \N__6893\,
            I => \N__6890\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__6890\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__6887\,
            I => \N__6884\
        );

    \I__612\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__6881\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__610\ : InMux
    port map (
            O => \N__6878\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__609\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6872\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__6872\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDCZ0Z3\
        );

    \I__607\ : InMux
    port map (
            O => \N__6869\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__606\ : InMux
    port map (
            O => \N__6866\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__605\ : InMux
    port map (
            O => \N__6863\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__604\ : InMux
    port map (
            O => \N__6860\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__603\ : InMux
    port map (
            O => \N__6857\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__6854\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2_cascade_\
        );

    \I__601\ : InMux
    port map (
            O => \N__6851\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__600\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__6845\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0\
        );

    \I__598\ : InMux
    port map (
            O => \N__6842\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__597\ : IoInMux
    port map (
            O => \N__6839\,
            I => \N__6836\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__595\ : IoSpan4Mux
    port map (
            O => \N__6833\,
            I => \N__6830\
        );

    \I__594\ : Odrv4
    port map (
            O => \N__6830\,
            I => \Clock12MHz_c\
        );

    \I__593\ : IoInMux
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__591\ : IoSpan4Mux
    port map (
            O => \N__6821\,
            I => \N__6818\
        );

    \I__590\ : IoSpan4Mux
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__589\ : IoSpan4Mux
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__588\ : Odrv4
    port map (
            O => \N__6812\,
            I => \Clock50MHz.PixelClock\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__586\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__6803\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__584\ : InMux
    port map (
            O => \N__6800\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_cry_7,
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_2_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un21_beamy_cry_8,
            carryinitout => \bfn_2_13_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_4_0_\
        );

    \IN_MUX_bfv_2_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_4_0_\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_4_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_7_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_3_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6827\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8462\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9116\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_4_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BAT_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7617\,
            in2 => \N__6809\,
            in3 => \N__6800\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI7BATZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVH1_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7541\,
            in2 => \N__7622\,
            in3 => \N__6866\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNI8FVHZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68E2_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7621\,
            in2 => \N__7727\,
            in3 => \N__6863\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJ68EZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIC29L5_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6956\,
            in1 => \N__7598\,
            in2 => \N__7709\,
            in3 => \N__6860\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQ2_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7688\,
            in2 => \_gnd_net_\,
            in3 => \N__6857\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2\,
            ltout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8LMQZ0Z2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRU85_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__6922\,
            in1 => \_gnd_net_\,
            in2 => \N__6854\,
            in3 => \_gnd_net_\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRRUZ0Z85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUUEM_0_8_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_RNIUUEM_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10239\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDC3_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6957\,
            in2 => \N__6896\,
            in3 => \N__6851\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNILPDCZ0Z3\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PU3_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6848\,
            in2 => \N__6962\,
            in3 => \N__6842\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIR5PUZ0Z3\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJ4_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6961\,
            in2 => \N__6941\,
            in3 => \N__6932\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNITBFJZ0Z4\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINP5QD_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7018\,
            in1 => \N__6929\,
            in2 => \N__6923\,
            in3 => \N__6908\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6905\,
            in2 => \_gnd_net_\,
            in3 => \N__6899\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4SZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9104\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10240\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10090\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8A6_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7013\,
            in2 => \N__6887\,
            in3 => \N__6878\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIDH8AZ0Z6\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RH9_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6875\,
            in2 => \N__7019\,
            in3 => \N__6869\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI31RHZ0Z9\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74A_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7017\,
            in2 => \N__7052\,
            in3 => \N__7043\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIAF74AZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIQGGSO_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7110\,
            in1 => \N__6995\,
            in2 => \N__7040\,
            in3 => \N__7031\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3E_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7028\,
            in2 => \_gnd_net_\,
            in3 => \N__7022\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIDPH3EZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUUEM_8_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__8315\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9261\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIRD4S5_0_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7012\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10946\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NE_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7070\,
            in2 => \N__7111\,
            in3 => \N__6989\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNI4J0NEZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATK_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7106\,
            in2 => \N__6986\,
            in3 => \N__6974\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNIBDATKZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4O_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6971\,
            in2 => \N__7112\,
            in3 => \N__6965\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI2VT4OZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7085\,
            in2 => \N__7121\,
            in3 => \N__7102\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CP_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7079\,
            in2 => \_gnd_net_\,
            in3 => \N__7073\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIEP3CPZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DSP2_0_8_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011011111001"
        )
    port map (
            in0 => \N__9295\,
            in1 => \N__8316\,
            in2 => \N__12112\,
            in3 => \N__7270\,
            lcout => \beamY_RNI9DSP2_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10104\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICLER6_8_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7163\,
            in1 => \N__7058\,
            in2 => \_gnd_net_\,
            in3 => \N__8306\,
            lcout => chary_if_generate_plus_mult1_un47_sum_axb4,
            ltout => \chary_if_generate_plus_mult1_un47_sum_axb4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKM9GC_9_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111010000"
        )
    port map (
            in0 => \N__12236\,
            in1 => \N__7269\,
            in2 => \N__7064\,
            in3 => \N__7157\,
            lcout => OPEN,
            ltout => \beamY_RNIKM9GCZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI42CCP_5_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7148\,
            in2 => \N__7061\,
            in3 => \N__8461\,
            lcout => chary_if_generate_plus_mult1_un47_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIM5433_8_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__12233\,
            in1 => \N__9298\,
            in2 => \N__7278\,
            in3 => \N__12059\,
            lcout => \beamY_RNIM5433Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI93821_9_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__9296\,
            in1 => \N__7795\,
            in2 => \_gnd_net_\,
            in3 => \N__9608\,
            lcout => \beamY_RNI93821Z0Z_9\,
            ltout => \beamY_RNI93821Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIM5433_0_8_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101101001"
        )
    port map (
            in0 => \N__12234\,
            in1 => \N__9297\,
            in2 => \N__7166\,
            in3 => \N__12058\,
            lcout => \beamY_RNIM5433_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIIR4K3_0_7_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8339\,
            in1 => \N__7286\,
            in2 => \_gnd_net_\,
            in3 => \N__8307\,
            lcout => \beamY_RNIIR4K3_0Z0Z_7\,
            ltout => \beamY_RNIIR4K3_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKM9GC_0_9_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__12235\,
            in1 => \N__7268\,
            in2 => \N__7151\,
            in3 => \N__7311\,
            lcout => \beamY_RNIKM9GC_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DSP2_8_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110110100"
        )
    port map (
            in0 => \N__12061\,
            in1 => \N__8311\,
            in2 => \N__7279\,
            in3 => \N__9344\,
            lcout => chary_if_generate_plus_mult1_un47_sum_axbxc5_2,
            ltout => \chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI41384_7_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001101001"
        )
    port map (
            in0 => \N__9482\,
            in1 => \N__8652\,
            in2 => \N__7142\,
            in3 => \N__12062\,
            lcout => OPEN,
            ltout => \beamY_RNI41384Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBDEO7_7_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__7139\,
            in1 => \N__12169\,
            in2 => \N__7130\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un54_sum_ac0_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIH5LL11_5_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100010000100"
        )
    port map (
            in0 => \N__8464\,
            in1 => \N__9105\,
            in2 => \N__7127\,
            in3 => \N__7189\,
            lcout => chary_if_generate_plus_mult1_un54_sum_ac0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIIGUB_4_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7903\,
            in1 => \N__7860\,
            in2 => \_gnd_net_\,
            in3 => \N__7834\,
            lcout => un8_beamylt9_0,
            ltout => \un8_beamylt9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI0A6L_7_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9672\,
            in1 => \N__7952\,
            in2 => \N__7124\,
            in3 => \N__7938\,
            lcout => un5_visibley_c6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIIQEC2_9_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__7274\,
            in1 => \N__8463\,
            in2 => \_gnd_net_\,
            in3 => \N__12244\,
            lcout => chary_if_generate_plus_mult1_un47_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIP8FF1_1_7_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101101001"
        )
    port map (
            in0 => \N__9481\,
            in1 => \N__8651\,
            in2 => \N__9353\,
            in3 => \N__12060\,
            lcout => \beamY_RNIP8FF1_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUFT79_9_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110000110110"
        )
    port map (
            in0 => \N__7280\,
            in1 => \N__7330\,
            in2 => \N__8488\,
            in3 => \N__12254\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb4_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2BHS32_9_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011000101101"
        )
    port map (
            in0 => \N__8481\,
            in1 => \N__7392\,
            in2 => \N__7775\,
            in3 => \N__7175\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axbxc5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBV5E51_0_8_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__7224\,
            in1 => \N__7326\,
            in2 => \N__7368\,
            in3 => \N__7203\,
            lcout => \beamY_RNIBV5E51_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBV5E51_8_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7204\,
            in1 => \N__7360\,
            in2 => \N__7334\,
            in3 => \N__7225\,
            lcout => OPEN,
            ltout => \beamY_RNIBV5E51Z0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI8QGGE2_8_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8270\,
            in2 => \N__7235\,
            in3 => \N__7232\,
            lcout => chary_if_generate_plus_mult1_un54_sum_axbxc5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIRV5601_8_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8269\,
            in1 => \N__8479\,
            in2 => \N__7205\,
            in3 => \N__7226\,
            lcout => chary_if_generate_plus_mult1_un54_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVADQV_8_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8263\,
            in1 => \N__7223\,
            in2 => \_gnd_net_\,
            in3 => \N__7199\,
            lcout => \beamY_RNIVADQVZ0Z_8\,
            ltout => \beamY_RNIVADQVZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2BHS32_0_9_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111100100110"
        )
    port map (
            in0 => \N__7771\,
            in1 => \N__8480\,
            in2 => \N__7178\,
            in3 => \N__7174\,
            lcout => chary_if_generate_plus_mult1_un54_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIV5SUC3_0_9_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__7332\,
            in1 => \N__7367\,
            in2 => \N__8571\,
            in3 => \N__7394\,
            lcout => OPEN,
            ltout => \beamY_RNIV5SUC3_0Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0N9QT8_9_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8740\,
            in2 => \N__7409\,
            in3 => \N__7295\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axbxc5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI3SC791_5_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9110\,
            in1 => \N__7390\,
            in2 => \N__7369\,
            in3 => \N__7331\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIURID92_5_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7391\,
            in1 => \N__9111\,
            in2 => \N__7406\,
            in3 => \N__8786\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb4_0,
            ltout => \chary_if_generate_plus_mult1_un61_sum_axb4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIEIALM5_4_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000001000"
        )
    port map (
            in0 => \N__10243\,
            in1 => \N__7503\,
            in2 => \N__7397\,
            in3 => \N__8556\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_7_d,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_13_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100111110000"
        )
    port map (
            in0 => \N__8557\,
            in1 => \N__8609\,
            in2 => \N__8807\,
            in3 => \N__9112\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIV5SUC3_9_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7393\,
            in1 => \N__8552\,
            in2 => \N__7370\,
            in3 => \N__7333\,
            lcout => \beamY_RNIV5SUC3Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIB6AOI5_5_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000011100"
        )
    port map (
            in0 => \N__8614\,
            in1 => \N__8806\,
            in2 => \N__9122\,
            in3 => \N__8579\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0,
            ltout => \chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ0797K_4_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__8521\,
            in1 => \N__9984\,
            in2 => \N__7289\,
            in3 => \N__9852\,
            lcout => \beamY_RNIJ0797KZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g1_0_0_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001101001"
        )
    port map (
            in0 => \N__9988\,
            in1 => \N__10260\,
            in2 => \N__7463\,
            in3 => \N__8524\,
            lcout => g1_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g1_1_0_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10259\,
            in1 => \N__10321\,
            in2 => \_gnd_net_\,
            in3 => \N__9987\,
            lcout => g1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGMN7D3_4_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__10253\,
            in1 => \N__7504\,
            in2 => \_gnd_net_\,
            in3 => \N__8580\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axb4_0,
            ltout => \chary_if_generate_plus_mult1_un68_sum_axb4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI96MFKN_4_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__8522\,
            in1 => \N__7441\,
            in2 => \N__7454\,
            in3 => \N__9985\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axb4_i,
            ltout => \chary_if_generate_plus_mult1_un68_sum_axb4_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g2_1_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__11377\,
            in1 => \N__11827\,
            in2 => \N__7451\,
            in3 => \N__7448\,
            lcout => g2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_4_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000100011110"
        )
    port map (
            in0 => \N__8523\,
            in1 => \N__7442\,
            in2 => \N__7433\,
            in3 => \N__9986\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axb4_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g2_0_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000000000"
        )
    port map (
            in0 => \N__11376\,
            in1 => \N__7424\,
            in2 => \N__11831\,
            in3 => \N__7418\,
            lcout => OPEN,
            ltout => \g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_7_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__8729\,
            in1 => \N__7529\,
            in2 => \N__7412\,
            in3 => \N__10322\,
            lcout => chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI074AD4_5_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7522\,
            in2 => \_gnd_net_\,
            in3 => \N__8578\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb4_i,
            ltout => \chary_if_generate_plus_mult1_un61_sum_axb4_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_2_0_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11823\,
            in1 => \N__8695\,
            in2 => \N__7532\,
            in3 => \N__10016\,
            lcout => \un114_pixel_6_1_5__g0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIRLTLI4_0_5_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111010100"
        )
    port map (
            in0 => \N__9120\,
            in1 => \N__8613\,
            in2 => \N__10261\,
            in3 => \N__8577\,
            lcout => chary_if_generate_plus_mult1_un61_sum_c4,
            ltout => \chary_if_generate_plus_mult1_un61_sum_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISDTA58_5_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__7523\,
            in1 => \_gnd_net_\,
            in2 => \N__7511\,
            in3 => \N__7508\,
            lcout => OPEN,
            ltout => \beamY_RNISDTA58Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0DLMCS_3_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__11822\,
            in1 => \N__11375\,
            in2 => \N__7487\,
            in3 => \N__7484\,
            lcout => chary_if_generate_plus_mult1_un75_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7592\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVL21_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7469\,
            in2 => \N__14251\,
            in3 => \N__7478\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNICVLZ0Z21\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1N21_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12102\,
            in2 => \N__14252\,
            in3 => \N__7475\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNID1NZ0Z21\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7472\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2B511_0_9_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12101\,
            lcout => \beamY_RNI2B511_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12255\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6U_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7583\,
            in2 => \N__14275\,
            in3 => \N__7577\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI6S6UZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEA1_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7574\,
            in2 => \N__14277\,
            in3 => \N__7568\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNILUEAZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HA1_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7565\,
            in2 => \N__14276\,
            in3 => \N__7559\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIN2HAZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7677\,
            in2 => \_gnd_net_\,
            in3 => \N__7556\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7550\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7553\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTEZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7549\,
            in2 => \_gnd_net_\,
            in3 => \N__7678\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_axb_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8482\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_4_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONL_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7784\,
            in2 => \N__7651\,
            in3 => \N__7535\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI4ONLZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVH1_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7646\,
            in2 => \N__7736\,
            in3 => \N__7718\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIEDVHZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8U1_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7715\,
            in2 => \N__7652\,
            in3 => \N__7700\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUH8UZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINI2Q2_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7616\,
            in1 => \N__7628\,
            in2 => \N__7697\,
            in3 => \N__7682\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7650\,
            in1 => \N__7679\,
            in2 => \N__7664\,
            in3 => \N__7655\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMRZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNIOTE9_0_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7642\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIMQMR_0_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7615\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9260\,
            in2 => \_gnd_net_\,
            in3 => \N__8318\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb3_i_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_axb3_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010010100"
        )
    port map (
            in0 => \N__12257\,
            in1 => \N__12154\,
            in2 => \N__8489\,
            in3 => \N__12082\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_axbZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12256\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIM5M02_9_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100110100110"
        )
    port map (
            in0 => \N__12259\,
            in1 => \N__9328\,
            in2 => \N__7802\,
            in3 => \N__9588\,
            lcout => chary_if_generate_plus_mult1_un47_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_8_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8141\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13139\,
            ce => \N__11545\,
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_6_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100111"
        )
    port map (
            in0 => \N__12084\,
            in1 => \N__12260\,
            in2 => \N__12173\,
            in3 => \N__8475\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_axb4_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010001001001"
        )
    port map (
            in0 => \N__12258\,
            in1 => \N__12158\,
            in2 => \N__8487\,
            in3 => \N__12083\,
            lcout => row_1_if_generate_plus_mult1_un61_sum_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIF0BK31_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__7757\,
            in1 => \N__10947\,
            in2 => \_gnd_net_\,
            in3 => \N__7748\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__10948\,
            in1 => \N__14278\,
            in2 => \_gnd_net_\,
            in3 => \N__11321\,
            lcout => \beamY_i_2\,
            ltout => \beamY_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_1_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010001000"
        )
    port map (
            in0 => \N__7756\,
            in1 => \N__7747\,
            in2 => \N__7739\,
            in3 => \N__10903\,
            lcout => \un114_pixel_6_1_5__chessboardpixel_un200_pixellto4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_3_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8051\,
            in2 => \_gnd_net_\,
            in3 => \N__11446\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13138\,
            ce => \N__11530\,
            sr => \_gnd_net_\
        );

    \beamY_fast_3_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8047\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11428\,
            lcout => \beamY_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13136\,
            ce => \N__11543\,
            sr => \_gnd_net_\
        );

    \beamY_fast_6_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7988\,
            lcout => \beamY_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13136\,
            ce => \N__11543\,
            sr => \_gnd_net_\
        );

    \beamY_fast_8_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8137\,
            lcout => \beamY_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13136\,
            ce => \N__11543\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7966\,
            in2 => \_gnd_net_\,
            in3 => \N__11427\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13136\,
            ce => \N__11543\,
            sr => \_gnd_net_\
        );

    \beamY_fast_7_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__11430\,
            in1 => \_gnd_net_\,
            in2 => \N__7970\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13136\,
            ce => \N__11543\,
            sr => \_gnd_net_\
        );

    \beamY_fast_4_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__8027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11429\,
            lcout => \beamY_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13136\,
            ce => \N__11543\,
            sr => \_gnd_net_\
        );

    \beamY_RNID2EU_6_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__9491\,
            in1 => \N__9411\,
            in2 => \_gnd_net_\,
            in3 => \N__7811\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIT5UF_4_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__7939\,
            in1 => \N__7918\,
            in2 => \N__7904\,
            in3 => \N__7833\,
            lcout => OPEN,
            ltout => \beamY_fast_RNIT5UFZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIKRSR_5_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100010"
        )
    port map (
            in0 => \N__7919\,
            in1 => \N__7940\,
            in2 => \N__7814\,
            in3 => \N__7861\,
            lcout => un5_visibley_ac0_7,
            ltout => \un5_visibley_ac0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICOMV_6_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010111"
        )
    port map (
            in0 => \N__9607\,
            in1 => \N__9412\,
            in2 => \N__7805\,
            in3 => \N__9492\,
            lcout => chary_if_generate_plus_mult1_un40_sum_axbxc5_i2_mux,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_5_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8006\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13134\,
            ce => \N__11555\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI6FUF_7_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7951\,
            in1 => \N__7937\,
            in2 => \N__7886\,
            in3 => \N__7917\,
            lcout => OPEN,
            ltout => \un5_visibley_ac0_11_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2B511_9_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9606\,
            in2 => \N__7907\,
            in3 => \N__7871\,
            lcout => chary_if_generate_plus_mult1_un33_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIT5UF_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7899\,
            in1 => \N__7859\,
            in2 => \N__7885\,
            in3 => \N__7832\,
            lcout => un5_visibley_c7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8065\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13135\,
            ce => \N__11544\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8026\,
            in2 => \_gnd_net_\,
            in3 => \N__11447\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13135\,
            ce => \N__11544\,
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un8_beamylto4_0_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7865\,
            in2 => \_gnd_net_\,
            in3 => \N__7835\,
            lcout => un5_visibley_c2,
            ltout => \un5_visibley_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISKOB_5_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__9798\,
            in1 => \N__9409\,
            in2 => \N__7838\,
            in3 => \N__9670\,
            lcout => un5_visibley_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_2_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8066\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13135\,
            ce => \N__11544\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7984\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13137\,
            ce => \N__11554\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8002\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13137\,
            ce => \N__11554\,
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15132\,
            in2 => \N__14939\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => un21_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_RNIAL73_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11378\,
            in2 => \_gnd_net_\,
            in3 => \N__8054\,
            lcout => \un21_beamy_cry_1_c_RNIALZ0Z73\,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => un21_beamy_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_2_c_RNICO83_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11810\,
            in2 => \_gnd_net_\,
            in3 => \N__8030\,
            lcout => \un21_beamy_cry_2_c_RNICOZ0Z83\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_3_c_RNIER93_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9839\,
            in2 => \_gnd_net_\,
            in3 => \N__8009\,
            lcout => \un21_beamy_cry_3_c_RNIERZ0Z93\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_4_c_RNIGUA3_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9671\,
            in2 => \_gnd_net_\,
            in3 => \N__7991\,
            lcout => \un21_beamy_cry_4_c_RNIGUAZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_5_c_RNII1C3_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9410\,
            in2 => \_gnd_net_\,
            in3 => \N__7973\,
            lcout => \un21_beamy_cry_5_c_RNII1CZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_6_c_RNIK4D3_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9510\,
            in2 => \_gnd_net_\,
            in3 => \N__7955\,
            lcout => \un21_beamy_cry_6_c_RNIK4DZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_7_c_RNIM7E3_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9340\,
            in2 => \_gnd_net_\,
            in3 => \N__8120\,
            lcout => \un21_beamy_cry_7_c_RNIM7EZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_9_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__9605\,
            in1 => \N__11453\,
            in2 => \_gnd_net_\,
            in3 => \N__8117\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13140\,
            ce => \N__11546\,
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14238\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9148\,
            lcout => if_generate_plus_mult1_un61_sum_axbxc5,
            ltout => \if_generate_plus_mult1_un61_sum_axbxc5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011001111001"
        )
    port map (
            in0 => \N__9097\,
            in1 => \N__8110\,
            in2 => \N__8114\,
            in3 => \N__8234\,
            lcout => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_7_0_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010110110010"
        )
    port map (
            in0 => \N__9096\,
            in1 => \N__10372\,
            in2 => \N__8111\,
            in3 => \N__8233\,
            lcout => row_1_if_generate_plus_mult1_un68_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_ac0_5_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100010000010"
        )
    port map (
            in0 => \N__10241\,
            in1 => \N__9149\,
            in2 => \N__14271\,
            in3 => \N__9095\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_ac0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_7_d_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__8089\,
            in1 => \N__8235\,
            in2 => \_gnd_net_\,
            in3 => \N__9072\,
            lcout => OPEN,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_ac0_7_dZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110101"
        )
    port map (
            in0 => \N__8246\,
            in1 => \N__10396\,
            in2 => \N__8096\,
            in3 => \N__8471\,
            lcout => row_1_if_generate_plus_mult1_un61_sum_c5,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m5_i_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__14272\,
            in1 => \_gnd_net_\,
            in2 => \N__8093\,
            in3 => \N__9075\,
            lcout => \row_1_if_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_0_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100111000011"
        )
    port map (
            in0 => \N__9073\,
            in1 => \N__8090\,
            in2 => \N__8078\,
            in3 => \N__8237\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_1_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011011101"
        )
    port map (
            in0 => \N__12271\,
            in1 => \N__12174\,
            in2 => \_gnd_net_\,
            in3 => \N__12108\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_ac0_7_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_m5x_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9074\,
            in1 => \N__14273\,
            in2 => \N__10262\,
            in3 => \N__9150\,
            lcout => row_1_if_i4_mux_i,
            ltout => \row_1_if_i4_mux_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011010001001"
        )
    port map (
            in0 => \N__10242\,
            in1 => \N__8185\,
            in2 => \N__8240\,
            in3 => \N__8236\,
            lcout => OPEN,
            ltout => \row_1_if_generate_plus_mult1_un75_sum_ac0_7_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_ac0_7_0_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__10094\,
            in1 => \N__8204\,
            in2 => \N__8198\,
            in3 => \N__8195\,
            lcout => row_1_if_generate_plus_mult1_un75_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10257\,
            in1 => \N__11008\,
            in2 => \N__10096\,
            in3 => \N__11049\,
            lcout => if_generate_plus_mult1_un75_sum_axbxc3,
            ltout => \if_generate_plus_mult1_un75_sum_axbxc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axb4_x0_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11050\,
            in1 => \N__8163\,
            in2 => \N__8189\,
            in3 => \N__11009\,
            lcout => if_generate_plus_mult1_un82_sum_axb4_x0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__14274\,
            in1 => \N__8186\,
            in2 => \_gnd_net_\,
            in3 => \N__9151\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\,
            ltout => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8164\,
            in1 => \N__8357\,
            in2 => \N__8171\,
            in3 => \N__11052\,
            lcout => if_generate_plus_mult1_un75_sum_axbxc5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axb4_x1_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11051\,
            in1 => \N__11010\,
            in2 => \N__8168\,
            in3 => \N__8147\,
            lcout => OPEN,
            ltout => \if_generate_plus_mult1_un82_sum_axb4_x1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axb4_ns_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8356\,
            in2 => \N__8348\,
            in3 => \N__8345\,
            lcout => row_1_if_generate_plus_mult1_un82_sum_axb4_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIP8FF1_0_7_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__9499\,
            in1 => \N__9335\,
            in2 => \N__8673\,
            in3 => \N__12103\,
            lcout => \beamY_RNIP8FF1_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un5_beamx_3_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9846\,
            in1 => \N__15170\,
            in2 => \_gnd_net_\,
            in3 => \N__9336\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__un5_beamxZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un5_beamx_5_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14921\,
            in1 => \N__9500\,
            in2 => \N__8327\,
            in3 => \N__9625\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__un5_beamxZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un5_beamx_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9176\,
            in1 => \N__11772\,
            in2 => \N__8324\,
            in3 => \N__11329\,
            lcout => un5_beamx_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_5_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__11328\,
            in1 => \N__9845\,
            in2 => \N__11809\,
            in3 => \N__9691\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un54_sum_axbxc5_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110110011011"
        )
    port map (
            in0 => \N__12270\,
            in1 => \N__12176\,
            in2 => \N__8486\,
            in3 => \N__12104\,
            lcout => if_generate_plus_mult1_un54_sum_axbxc5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIP8FF1_7_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101101"
        )
    port map (
            in0 => \N__9522\,
            in1 => \N__9346\,
            in2 => \N__8675\,
            in3 => \N__12091\,
            lcout => OPEN,
            ltout => \beamY_RNIP8FF1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIIR4K3_7_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8630\,
            in2 => \N__8321\,
            in3 => \N__8317\,
            lcout => chary_if_generate_plus_mult1_un40_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIP8FF1_2_7_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110111"
        )
    port map (
            in0 => \N__9521\,
            in1 => \N__9345\,
            in2 => \N__8674\,
            in3 => \N__12090\,
            lcout => \beamY_RNIP8FF1_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_0_3_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11781\,
            in2 => \_gnd_net_\,
            in3 => \N__11366\,
            lcout => OPEN,
            ltout => \un4_beamylt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_beamylto6_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9847\,
            in1 => \N__9426\,
            in2 => \N__8624\,
            in3 => \N__9692\,
            lcout => un4_beamylt8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un8_beamylto9_0_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9350\,
            in1 => \N__9523\,
            in2 => \_gnd_net_\,
            in3 => \N__9609\,
            lcout => \un114_pixel_6_1_5__un8_beamylto9Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIRLTLI4_5_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8621\,
            in1 => \N__9109\,
            in2 => \N__10249\,
            in3 => \N__8582\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c5_0_i4_mux_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIB6AOI5_0_5_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000011100"
        )
    port map (
            in0 => \N__8620\,
            in1 => \N__8808\,
            in2 => \N__9121\,
            in3 => \N__8581\,
            lcout => OPEN,
            ltout => \beamY_RNIB6AOI5_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPOKD9B_5_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8528\,
            in3 => \N__8525\,
            lcout => chary_if_generate_plus_mult1_un61_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISKOB_0_5_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010010011"
        )
    port map (
            in0 => \N__8501\,
            in1 => \N__9413\,
            in2 => \N__9853\,
            in3 => \N__9673\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI3GESM7_4_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000101010"
        )
    port map (
            in0 => \N__8764\,
            in1 => \N__8809\,
            in2 => \N__10238\,
            in3 => \N__8752\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c5_0,
            ltout => \chary_if_generate_plus_mult1_un68_sum_c5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_11_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__8825\,
            in1 => \N__11815\,
            in2 => \N__8816\,
            in3 => \N__11593\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un1_sum_axbxc3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_0_5_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110110111100"
        )
    port map (
            in0 => \N__8714\,
            in1 => \N__14920\,
            in2 => \N__8813\,
            in3 => \N__11367\,
            lcout => \un114_pixel_6_1_5__font_un126_pixel_m_4_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNILT8E7K_3_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111010100"
        )
    port map (
            in0 => \N__10198\,
            in1 => \N__10301\,
            in2 => \N__10105\,
            in3 => \N__10020\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI3GESM7_0_4_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110001001100"
        )
    port map (
            in0 => \N__8810\,
            in1 => \N__8765\,
            in2 => \N__10258\,
            in3 => \N__8753\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c5_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_17_1_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111101010"
        )
    port map (
            in0 => \N__10853\,
            in1 => \N__8681\,
            in2 => \N__10106\,
            in3 => \N__11677\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__g0_17Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_17_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9717\,
            in1 => \N__11592\,
            in2 => \N__8717\,
            in3 => \N__9746\,
            lcout => chary_if_generate_plus_mult1_un75_sum_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKC087T_5_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__8708\,
            in1 => \N__10310\,
            in2 => \N__8699\,
            in3 => \N__10021\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axbxc5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4VNB7K_0_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__10022\,
            in1 => \_gnd_net_\,
            in2 => \N__10320\,
            in3 => \N__10237\,
            lcout => g1_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15279\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5J6_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8860\,
            in2 => \N__10352\,
            in3 => \N__8873\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8E5JZ0Z6\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQ9_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9929\,
            in2 => \N__9896\,
            in3 => \N__8870\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIEEGQZ0Z9\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI17AMN_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8923\,
            in1 => \N__8861\,
            in2 => \N__9920\,
            in3 => \N__8867\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9908\,
            in2 => \_gnd_net_\,
            in3 => \N__8864\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BCZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_0_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9891\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16131\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_5_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGC_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8903\,
            in2 => \N__8897\,
            in3 => \N__8852\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIGSPGCZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1J_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8849\,
            in2 => \N__8924\,
            in3 => \N__8843\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNI0CU1JZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8831\,
            in2 => \N__8840\,
            in3 => \N__8919\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_invZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPN_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8933\,
            in2 => \_gnd_net_\,
            in3 => \N__8927\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIEVUPNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNID96BC_0_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8918\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_1_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15280\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10487\,
            in2 => \N__14497\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10518\,
            in2 => \_gnd_net_\,
            in3 => \N__8888\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__13145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10736\,
            in2 => \_gnd_net_\,
            in3 => \N__8885\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__13145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11509\,
            in1 => \N__10772\,
            in2 => \_gnd_net_\,
            in3 => \N__8882\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__13145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10686\,
            in2 => \_gnd_net_\,
            in3 => \N__8879\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__13145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10564\,
            in2 => \_gnd_net_\,
            in3 => \N__8876\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__13145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11171\,
            in2 => \_gnd_net_\,
            in3 => \N__8972\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__13145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10634\,
            in2 => \_gnd_net_\,
            in3 => \N__8969\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__13145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10600\,
            in2 => \_gnd_net_\,
            in3 => \N__8966\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__13142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11138\,
            in1 => \N__11508\,
            in2 => \_gnd_net_\,
            in3 => \N__8963\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_row_1_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101000101"
        )
    port map (
            in0 => \N__8960\,
            in1 => \N__11808\,
            in2 => \N__10095\,
            in3 => \N__11365\,
            lcout => \un114_pixel_6_1_5__un4_rowZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un3_beamx_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__11190\,
            in1 => \N__11170\,
            in2 => \N__10690\,
            in3 => \N__10358\,
            lcout => un3_beamx_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un15_beamy_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__8954\,
            in1 => \N__8945\,
            in2 => \N__11139\,
            in3 => \N__9174\,
            lcout => \un114_pixel_6_1_5__un15_beamyZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un1_beamxlto6_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10739\,
            in1 => \N__10694\,
            in2 => \N__10778\,
            in3 => \N__10568\,
            lcout => un1_beamxlt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un1_beamylto9_0_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9851\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11796\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__un1_beamylto9Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un1_beamylto9_3_0_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__11330\,
            in1 => \N__14922\,
            in2 => \N__9215\,
            in3 => \N__9501\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__un1_beamylto9_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__9175\,
            in1 => \N__9349\,
            in2 => \N__9212\,
            in3 => \N__9626\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un3_beamx_2_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10598\,
            in2 => \_gnd_net_\,
            in3 => \N__10637\,
            lcout => un1_beamx_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_20_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__9624\,
            in1 => \N__9525\,
            in2 => \N__8987\,
            in3 => \N__9348\,
            lcout => un4_beamy_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un5_beamx_4_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9425\,
            in2 => \_gnd_net_\,
            in3 => \N__9688\,
            lcout => un8_beamy_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11780\,
            in2 => \_gnd_net_\,
            in3 => \N__11368\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum,
            ltout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_1_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011101001101"
        )
    port map (
            in0 => \N__10212\,
            in1 => \N__11017\,
            in2 => \N__9161\,
            in3 => \N__11059\,
            lcout => OPEN,
            ltout => \row_1_if_generate_plus_mult1_un82_sum_axbxc5_3Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_3_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__14279\,
            in1 => \N__9158\,
            in2 => \N__9125\,
            in3 => \N__9062\,
            lcout => \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_beamylto9_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__9623\,
            in1 => \N__9524\,
            in2 => \N__8986\,
            in3 => \N__9347\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_1_4_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9689\,
            in1 => \N__9526\,
            in2 => \N__9431\,
            in3 => \N__11794\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__g0_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_0_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100000000"
        )
    port map (
            in0 => \N__9616\,
            in1 => \N__9224\,
            in2 => \N__9695\,
            in3 => \N__14499\,
            lcout => \un114_pixel_6_1_5__g0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_0_4_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9690\,
            in1 => \N__9351\,
            in2 => \N__9854\,
            in3 => \N__9615\,
            lcout => \un114_pixel_6_1_5__g0_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_0_3_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__11795\,
            in1 => \_gnd_net_\,
            in2 => \N__9530\,
            in3 => \N__9430\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__g0_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_8_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__9368\,
            in1 => \N__14854\,
            in2 => \N__9359\,
            in3 => \N__11374\,
            lcout => un1_beamy_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g2_0_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__11332\,
            in1 => \N__11782\,
            in2 => \_gnd_net_\,
            in3 => \N__11672\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__g2_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJH2N2P_0_3_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111101010"
        )
    port map (
            in0 => \N__10854\,
            in1 => \N__9860\,
            in2 => \N__9356\,
            in3 => \N__9767\,
            lcout => \N_80_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ3MRIJ1_3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000011110"
        )
    port map (
            in0 => \N__9953\,
            in1 => \N__10855\,
            in2 => \N__11811\,
            in3 => \N__11673\,
            lcout => m511_0_o2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_0_1_1_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__9844\,
            in1 => \N__11333\,
            in2 => \N__14898\,
            in3 => \N__9352\,
            lcout => \un114_pixel_6_1_5__g0_0_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4VNB7K_1_4_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__10199\,
            in1 => \N__10305\,
            in2 => \_gnd_net_\,
            in3 => \N__10017\,
            lcout => g1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_4_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__9843\,
            in1 => \N__11776\,
            in2 => \_gnd_net_\,
            in3 => \N__11331\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum,
            ltout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4VNB7K_4_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10306\,
            in2 => \N__9770\,
            in3 => \N__10018\,
            lcout => g1_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIITKSF53_3_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11589\,
            in1 => \N__9713\,
            in2 => \N__11671\,
            in3 => \N__9747\,
            lcout => m511_0_x2_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ3MRIJ1_0_3_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101011010"
        )
    port map (
            in0 => \N__10861\,
            in1 => \N__11658\,
            in2 => \N__11828\,
            in3 => \N__9952\,
            lcout => \G_7_0_m2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1KDQIJ1_3_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111101110"
        )
    port map (
            in0 => \N__9951\,
            in1 => \N__10860\,
            in2 => \_gnd_net_\,
            in3 => \N__11659\,
            lcout => OPEN,
            ltout => \G_7_0_m2_1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIABC7E1_3_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9749\,
            in1 => \N__9722\,
            in2 => \N__9761\,
            in3 => \N__11590\,
            lcout => OPEN,
            ltout => \G_7_0_m2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGABC8I2_2_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000100100"
        )
    port map (
            in0 => \N__11591\,
            in1 => \N__11380\,
            in2 => \N__9758\,
            in3 => \N__9755\,
            lcout => \G_7_0_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJH2N2P_3_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9748\,
            in1 => \N__11657\,
            in2 => \N__9721\,
            in3 => \N__9935\,
            lcout => \beamY_RNIJH2N2PZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNILT8E7K_0_3_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000010010000"
        )
    port map (
            in0 => \N__10295\,
            in1 => \N__10211\,
            in2 => \N__10097\,
            in3 => \N__10019\,
            lcout => chary_if_generate_plus_mult1_un68_sum_ac0_5,
            ltout => \chary_if_generate_plus_mult1_un68_sum_ac0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIL0E2QG2_3_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010110111010"
        )
    port map (
            in0 => \N__10859\,
            in1 => \N__11653\,
            in2 => \N__9938\,
            in3 => \N__11588\,
            lcout => \beamY_RNIL0E2QG2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14334\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02D93_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9868\,
            in2 => \N__9878\,
            in3 => \N__9923\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI02DZ0Z93\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVP4_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11878\,
            in2 => \N__11204\,
            in3 => \N__9911\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FVPZ0Z4\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIUPOTB_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9895\,
            in1 => \N__9869\,
            in2 => \N__11903\,
            in3 => \N__9902\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11O36_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11891\,
            in2 => \_gnd_net_\,
            in3 => \N__9899\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI11OZ0Z36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13678\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_0_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11877\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14335\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14476\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_5_0_\,
            carryout => un5_visiblex_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_RNIHKT1_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10489\,
            in3 => \N__10343\,
            lcout => charx_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_0,
            carryout => un5_visiblex_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10519\,
            in3 => \N__10340\,
            lcout => charx_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_1,
            carryout => un5_visiblex_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14236\,
            in2 => \N__10737\,
            in3 => \N__10337\,
            lcout => chessboardpixel_un152_pixel_24,
            ltout => OPEN,
            carryin => un5_visiblex_cry_2,
            carryout => un5_visiblex_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10773\,
            in3 => \N__10334\,
            lcout => charx_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_3,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10687\,
            in3 => \N__10331\,
            lcout => charx_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14237\,
            in2 => \N__10565\,
            in3 => \N__10328\,
            lcout => charx_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11162\,
            in2 => \_gnd_net_\,
            in3 => \N__10325\,
            lcout => charx_if_generate_plus_mult1_un33_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14266\,
            in2 => \N__10635\,
            in3 => \N__10412\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10594\,
            in2 => \_gnd_net_\,
            in3 => \N__10409\,
            lcout => \CO3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__14475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10488\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_1_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100010101"
        )
    port map (
            in0 => \N__10406\,
            in1 => \N__10810\,
            in2 => \N__16325\,
            in3 => \N__16135\,
            lcout => \un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14474\,
            in2 => \_gnd_net_\,
            in3 => \N__11507\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_row_5_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10400\,
            in1 => \N__10379\,
            in2 => \N__11999\,
            in3 => \N__12362\,
            lcout => \un114_pixel_6_1_5__un4_rowZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un3_beamx_5_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10771\,
            in1 => \N__10517\,
            in2 => \N__11140\,
            in3 => \N__10486\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__un3_beamxZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un3_beamx_7_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10563\,
            in1 => \N__10735\,
            in2 => \N__10361\,
            in3 => \N__14500\,
            lcout => \un114_pixel_6_1_5__un3_beamxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g3_0_1_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10599\,
            in2 => \_gnd_net_\,
            in3 => \N__10633\,
            lcout => \un114_pixel_6_1_5__g3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__chessboardpixel_un174_pixellto10_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001010010010"
        )
    port map (
            in0 => \N__10820\,
            in1 => \N__10814\,
            in2 => \N__10799\,
            in3 => \N__16145\,
            lcout => chessboardpixel_un174_pixel_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un13_beamylto7_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__11173\,
            in1 => \N__10689\,
            in2 => \N__10703\,
            in3 => \N__10567\,
            lcout => un13_beamylt10_0,
            ltout => \un13_beamylt10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un15_beamy_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100000000"
        )
    port map (
            in0 => \N__11191\,
            in1 => \N__10787\,
            in2 => \N__10781\,
            in3 => \N__10444\,
            lcout => un15_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un13_beamylto5_1_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__10774\,
            in1 => \N__10738\,
            in2 => \N__10454\,
            in3 => \N__14477\,
            lcout => un18_beamylt5_0,
            ltout => \un18_beamylt5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un15_beamy_1_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__10688\,
            in1 => \N__10529\,
            in2 => \N__10646\,
            in3 => \N__10643\,
            lcout => \un114_pixel_6_1_5__un15_beamyZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un18_beamylto9_2_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11172\,
            in1 => \N__10636\,
            in2 => \N__10601\,
            in3 => \N__10566\,
            lcout => \un114_pixel_6_1_5__un18_beamylto9Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un13_beamylto2_0_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10523\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10490\,
            lcout => \un114_pixel_6_1_5__un13_beamylto2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_19_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__10445\,
            in1 => \N__10436\,
            in2 => \N__10430\,
            in3 => \N__10418\,
            lcout => \un114_pixel_6_1_5__g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__11192\,
            in1 => \N__11174\,
            in2 => \N__11141\,
            in3 => \N__11108\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13144\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_row_7_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__11069\,
            in1 => \N__11060\,
            in2 => \N__11024\,
            in3 => \N__12434\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__un4_rowZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_row_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__10985\,
            in1 => \N__10973\,
            in2 => \N__10967\,
            in3 => \N__10964\,
            lcout => un4_row,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__chessboardpixel_un200_pixellto4_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__10955\,
            in1 => \N__10928\,
            in2 => \N__14905\,
            in3 => \N__10915\,
            lcout => OPEN,
            ltout => \chessboardpixel_un200_pixellt10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__chessboardpixel_un200_pixellto10_1_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001001"
        )
    port map (
            in0 => \N__10916\,
            in1 => \N__10892\,
            in2 => \N__10880\,
            in3 => \N__10877\,
            lcout => chessboardpixel_un200_pixel_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001101100"
        )
    port map (
            in0 => \N__11542\,
            in1 => \N__14855\,
            in2 => \N__15143\,
            in3 => \N__11448\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_1_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__11603\,
            in1 => \N__11615\,
            in2 => \N__11830\,
            in3 => \N__10865\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un1_sum_axbxc3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_0_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101010011110"
        )
    port map (
            in0 => \N__14847\,
            in1 => \N__11370\,
            in2 => \N__10823\,
            in3 => \N__11216\,
            lcout => \un114_pixel_6_1_5__font_un126_pixel_m_4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__11369\,
            in1 => \N__11837\,
            in2 => \N__11829\,
            in3 => \N__11678\,
            lcout => g2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_12_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12536\,
            in1 => \N__15107\,
            in2 => \_gnd_net_\,
            in3 => \N__13248\,
            lcout => \N_357_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPG1SS93_2_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011010010000"
        )
    port map (
            in0 => \N__11609\,
            in1 => \N__11602\,
            in2 => \N__11381\,
            in3 => \N__11561\,
            lcout => \beamY_RNIPG1SS93Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_i_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16439\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__15052\,
            in1 => \N__11553\,
            in2 => \_gnd_net_\,
            in3 => \N__11449\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_6_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__11379\,
            in1 => \N__11225\,
            in2 => \_gnd_net_\,
            in3 => \N__11215\,
            lcout => font_un28_pixel_0_0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13693\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_3_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILI1_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11854\,
            in2 => \N__11864\,
            in3 => \N__11195\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI1ILIZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLI2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12629\,
            in2 => \N__12596\,
            in3 => \N__11894\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIOPLIZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIP5RO5_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11879\,
            in1 => \N__11855\,
            in2 => \N__12620\,
            in3 => \N__11885\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FS2_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12608\,
            in2 => \_gnd_net_\,
            in3 => \N__11882\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNIU5FSZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_1_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13614\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_0_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12591\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14329\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_m_2_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__12713\,
            in1 => \N__13945\,
            in2 => \N__11942\,
            in3 => \N__11846\,
            lcout => if_generate_plus_mult1_un47_sum_m_2,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_1,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11933\,
            in2 => \N__12293\,
            in3 => \N__11843\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_3,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_2,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13946\,
            in2 => \N__12284\,
            in3 => \N__11840\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_4,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_3,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__13947\,
            in1 => \N__13609\,
            in2 => \N__13685\,
            in3 => \N__11948\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_5,
            ltout => \column_1_if_generate_plus_mult1_un47_sum1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_N_571_i_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12766\,
            in2 => \N__11945\,
            in3 => \N__13948\,
            lcout => \N_571_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_3_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13667\,
            lcout => un5_visiblex_i_0_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_3_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__13888\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un26_sum_axb_3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111000011"
        )
    port map (
            in0 => \N__12692\,
            in1 => \N__11974\,
            in2 => \N__11927\,
            in3 => \N__13893\,
            lcout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_m_5_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__13891\,
            in1 => \_gnd_net_\,
            in2 => \N__12748\,
            in3 => \N__12765\,
            lcout => if_generate_plus_mult1_un47_sum_m_5,
            ltout => \if_generate_plus_mult1_un47_sum_m_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110100101"
        )
    port map (
            in0 => \N__11915\,
            in1 => \N__12701\,
            in2 => \N__11909\,
            in3 => \N__13892\,
            lcout => OPEN,
            ltout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11906\,
            in3 => \N__12396\,
            lcout => if_generate_plus_mult1_un54_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_2_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13887\,
            lcout => \un5_visiblex_cry_8_c_RNI1D62Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m15_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__13889\,
            in1 => \N__13671\,
            in2 => \_gnd_net_\,
            in3 => \N__13591\,
            lcout => \N_11_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100110011"
        )
    port map (
            in0 => \N__13592\,
            in1 => \N__13552\,
            in2 => \N__13686\,
            in3 => \N__13890\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_m_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14330\,
            in2 => \N__14345\,
            in3 => \N__13886\,
            lcout => if_generate_plus_mult1_un47_sum_m_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_1_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13666\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_row_2_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__12275\,
            in1 => \N__12175\,
            in2 => \N__12731\,
            in3 => \N__12113\,
            lcout => \un114_pixel_6_1_5__un4_rowZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13918\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un26_sum_s_2_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15285\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12403\,
            in2 => \N__11990\,
            in3 => \N__11981\,
            lcout => if_generate_plus_mult1_un54_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11978\,
            in2 => \N__11963\,
            in3 => \N__11951\,
            lcout => if_generate_plus_mult1_un54_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12360\,
            in1 => \N__12416\,
            in2 => \N__12407\,
            in3 => \N__12383\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12380\,
            in2 => \_gnd_net_\,
            in3 => \N__12371\,
            lcout => if_generate_plus_mult1_un54_sum_s_5,
            ltout => \if_generate_plus_mult1_un54_sum_s_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12368\,
            in3 => \_gnd_net_\,
            lcout => column_1_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16156\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12331\,
            in2 => \N__12302\,
            in3 => \N__12365\,
            lcout => if_generate_plus_mult1_un61_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12361\,
            in2 => \N__12344\,
            in3 => \N__12335\,
            lcout => if_generate_plus_mult1_un61_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15385\,
            in1 => \N__12332\,
            in2 => \N__12323\,
            in3 => \N__12314\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12311\,
            in2 => \_gnd_net_\,
            in3 => \N__12305\,
            lcout => un5_rowlto3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_N_562_i_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15286\,
            lcout => \N_562_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__Pixel_3_sqmuxa_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001000000"
        )
    port map (
            in0 => \N__13039\,
            in1 => \N__12449\,
            in2 => \N__12892\,
            in3 => \N__12440\,
            lcout => \Pixel_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_rowlto3_sbtinv_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15383\,
            lcout => un5_rowlto3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_i_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16157\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_row_7_1_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__15685\,
            in1 => \N__16014\,
            in2 => \_gnd_net_\,
            in3 => \N__15384\,
            lcout => \un114_pixel_6_1_5__un4_row_7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI59CM492_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110011"
        )
    port map (
            in0 => \N__12428\,
            in1 => \N__16017\,
            in2 => \N__15233\,
            in3 => \N__13380\,
            lcout => OPEN,
            ltout => \N_18_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6M26DQ1_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__14848\,
            in1 => \_gnd_net_\,
            in2 => \N__12422\,
            in3 => \N__12461\,
            lcout => \N_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7LRQVE2_0_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101110111"
        )
    port map (
            in0 => \N__13097\,
            in1 => \N__16016\,
            in2 => \N__15162\,
            in3 => \N__13379\,
            lcout => OPEN,
            ltout => \N_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQVAMG32_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__14849\,
            in1 => \N__12479\,
            in2 => \N__12419\,
            in3 => \_gnd_net_\,
            lcout => \N_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_9_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001011111"
        )
    port map (
            in0 => \N__15862\,
            in1 => \N__14729\,
            in2 => \N__14929\,
            in3 => \N__16018\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__un116_pixel_3_1_0_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110100100100"
        )
    port map (
            in0 => \N__14850\,
            in1 => \N__12494\,
            in2 => \N__12482\,
            in3 => \N__13253\,
            lcout => \N_342_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISS6QGK3_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100001111"
        )
    port map (
            in0 => \N__12518\,
            in1 => \N__15106\,
            in2 => \N__12503\,
            in3 => \N__13374\,
            lcout => \N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m24_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15857\,
            in1 => \N__15665\,
            in2 => \_gnd_net_\,
            in3 => \N__16009\,
            lcout => column_0111_0,
            ltout => \column_0111_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI05CI5A3_0_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14382\,
            in2 => \N__12473\,
            in3 => \N__15101\,
            lcout => OPEN,
            ltout => \beamY_RNI05CI5A3_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBABJS01_1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__15102\,
            in1 => \N__14935\,
            in2 => \N__12470\,
            in3 => \N__12566\,
            lcout => OPEN,
            ltout => \beamY_RNIBABJS01Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__font_un126_pixel_2_am_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12644\,
            in2 => \N__12467\,
            in3 => \N__13373\,
            lcout => font_un126_pixel_2_am,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2QTJEJ1_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010010001"
        )
    port map (
            in0 => \N__15858\,
            in1 => \N__15666\,
            in2 => \N__15145\,
            in3 => \N__16010\,
            lcout => OPEN,
            ltout => \N_21_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIAVDE8H3_0_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15200\,
            in2 => \N__12464\,
            in3 => \N__13372\,
            lcout => \N_22_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNINIKJ5A3_1_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010111110"
        )
    port map (
            in0 => \N__14383\,
            in1 => \N__14934\,
            in2 => \N__15144\,
            in3 => \N__12455\,
            lcout => \beamY_RNINIKJ5A3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_3_bm_6_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011101000111"
        )
    port map (
            in0 => \N__15662\,
            in1 => \N__16048\,
            in2 => \N__15854\,
            in3 => \N__15481\,
            lcout => OPEN,
            ltout => \un116_pixel_3_bmZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISJITRQ2_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001110111"
        )
    port map (
            in0 => \N__14936\,
            in1 => \N__12542\,
            in2 => \N__12524\,
            in3 => \N__12509\,
            lcout => OPEN,
            ltout => \beamY_RNISJITRQ2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJDHE4C2_1_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__12548\,
            in1 => \_gnd_net_\,
            in2 => \N__12521\,
            in3 => \N__13371\,
            lcout => \beamY_RNIJDHE4C2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \m11_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110000000000"
        )
    port map (
            in0 => \N__15479\,
            in1 => \N__15806\,
            in2 => \N__16083\,
            in3 => \N__15663\,
            lcout => \N_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un114_pixel_3_i_m2_6_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011010011110"
        )
    port map (
            in0 => \N__15660\,
            in1 => \N__16038\,
            in2 => \N__15853\,
            in3 => \N__15477\,
            lcout => \un114_pixel_7_1_7__N_11_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m26_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__15478\,
            in1 => \N__15799\,
            in2 => \N__16082\,
            in3 => \N__15661\,
            lcout => OPEN,
            ltout => \N_248_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9GDVDD3_1_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__14873\,
            in1 => \N__15037\,
            in2 => \N__12512\,
            in3 => \N__13247\,
            lcout => un116_pixel_3_ns_1_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \m8_e_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100000000"
        )
    port map (
            in0 => \N__15480\,
            in1 => \N__15807\,
            in2 => \N__16084\,
            in3 => \N__15664\,
            lcout => \N_25_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__column_0001_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__16051\,
            in1 => \N__15655\,
            in2 => \N__15856\,
            in3 => \N__15471\,
            lcout => column_0001_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un114_pixel_3_i_a3_7_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__15656\,
            in1 => \N__15813\,
            in2 => \_gnd_net_\,
            in3 => \N__16053\,
            lcout => OPEN,
            ltout => \un114_pixel_3_i_a3_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI05CI5A3_0_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15036\,
            in2 => \N__12569\,
            in3 => \N__12562\,
            lcout => \beamY_RNI05CI5A3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2QTJEJ1_0_0_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010010001"
        )
    port map (
            in0 => \N__15653\,
            in1 => \N__15811\,
            in2 => \N__15097\,
            in3 => \N__16052\,
            lcout => OPEN,
            ltout => \un116_pixel_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDVSK5A3_1_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000110110"
        )
    port map (
            in0 => \N__14908\,
            in1 => \N__15035\,
            in2 => \N__12551\,
            in3 => \N__14380\,
            lcout => \beamY_RNIDVSK5A3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m12_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001000100"
        )
    port map (
            in0 => \N__16050\,
            in1 => \N__15654\,
            in2 => \N__15855\,
            in3 => \N__15470\,
            lcout => \N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_15_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011000000"
        )
    port map (
            in0 => \N__15469\,
            in1 => \N__15812\,
            in2 => \N__15684\,
            in3 => \N__16049\,
            lcout => \un114_pixel_0_1__N_6_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_4_bm_1_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011010111110"
        )
    port map (
            in0 => \N__16080\,
            in1 => \N__15594\,
            in2 => \N__15864\,
            in3 => \N__15473\,
            lcout => \un116_pixel_4_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_1_am_1_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010011111110111"
        )
    port map (
            in0 => \N__16079\,
            in1 => \N__14723\,
            in2 => \N__15863\,
            in3 => \N__15593\,
            lcout => OPEN,
            ltout => \un116_pixel_1_amZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUEM1HF2_1_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__14906\,
            in1 => \N__15000\,
            in2 => \N__12527\,
            in3 => \N__12635\,
            lcout => un116_pixel_3_ns_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_i_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16343\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_4_am_1_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100110011"
        )
    port map (
            in0 => \N__15474\,
            in1 => \N__15835\,
            in2 => \N__15659\,
            in3 => \N__16081\,
            lcout => OPEN,
            ltout => \un116_pixel_4_amZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHIRVUS1_1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__14907\,
            in1 => \N__12659\,
            in2 => \N__12653\,
            in3 => \N__12650\,
            lcout => \beamY_RNIHIRVUS1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_1_bm_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000011"
        )
    port map (
            in0 => \N__15472\,
            in1 => \N__15828\,
            in2 => \N__15658\,
            in3 => \N__16078\,
            lcout => \un116_pixel_1_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13613\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILF421_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12577\,
            in2 => \N__12722\,
            in3 => \N__12623\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNILFZ0Z421\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPB1_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13736\,
            in2 => \N__13757\,
            in3 => \N__12611\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNINJPBZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIKJPN2_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12595\,
            in1 => \N__12578\,
            in2 => \N__13724\,
            in3 => \N__12602\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTB1_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__13756\,
            in1 => \N__13712\,
            in2 => \_gnd_net_\,
            in3 => \N__12599\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIRRTBZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_0_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13752\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13956\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14350\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12674\,
            in2 => \N__12776\,
            in3 => \N__12704\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_2,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_1,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12680\,
            in2 => \N__12785\,
            in3 => \N__12695\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_3,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_2,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13742\,
            in2 => \N__12668\,
            in3 => \N__12686\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_4,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_3,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13955\,
            in2 => \_gnd_net_\,
            in3 => \N__12683\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__13953\,
            in1 => \_gnd_net_\,
            in2 => \N__13550\,
            in3 => \_gnd_net_\,
            lcout => if_generate_plus_mult1_un47_sum_0_cry_3_ma,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \N__13694\,
            in1 => \N__13535\,
            in2 => \_gnd_net_\,
            in3 => \N__13952\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__N_200_0_i_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__13954\,
            in1 => \_gnd_net_\,
            in2 => \N__13551\,
            in3 => \_gnd_net_\,
            lcout => \N_200_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13616\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12815\,
            in3 => \N__12806\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIH538_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14184\,
            in2 => \N__12803\,
            in3 => \N__12794\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNIHZ0Z538\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_LUT4_0_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13961\,
            in3 => \N__12791\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_LUT4_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12788\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__13684\,
            in1 => \N__13507\,
            in2 => \N__13553\,
            in3 => \N__13960\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_2_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13683\,
            lcout => un5_visiblex_i_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un4_row_0_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__13546\,
            in1 => \N__12767\,
            in2 => \N__12749\,
            in3 => \N__13959\,
            lcout => \un114_pixel_6_1_5__un4_rowZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13605\,
            lcout => un5_visiblex_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16446\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_5_bm_6_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100111100"
        )
    port map (
            in0 => \N__15411\,
            in1 => \N__15869\,
            in2 => \N__16086\,
            in3 => \N__15682\,
            lcout => \un116_pixel_5_bmZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_5_am_6_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011011011110"
        )
    port map (
            in0 => \N__15683\,
            in1 => \N__16070\,
            in2 => \N__15875\,
            in3 => \N__15412\,
            lcout => OPEN,
            ltout => \un116_pixel_5_amZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII25UDD3_0_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15166\,
            in2 => \N__12902\,
            in3 => \N__12899\,
            lcout => \beamY_RNII25UDD3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__font_un126_pixel_m_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__12893\,
            in1 => \N__14545\,
            in2 => \_gnd_net_\,
            in3 => \N__13387\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__font_un126_pixel_mZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_0_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__12872\,
            in1 => \N__14537\,
            in2 => \N__12860\,
            in3 => \N__14582\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__g0_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12857\,
            in2 => \N__12845\,
            in3 => \N__13046\,
            lcout => \Pixel_1_r_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g1_0_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__13388\,
            in1 => \_gnd_net_\,
            in2 => \N__14549\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \un114_pixel_6_1_5__g1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_16_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12842\,
            in1 => \N__12830\,
            in2 => \N__12818\,
            in3 => \N__13045\,
            lcout => \un114_pixel_6_1_5__font_un126_pixel_m_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIP6FOQ73_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13028\,
            in1 => \N__13016\,
            in2 => \_gnd_net_\,
            in3 => \N__13010\,
            lcout => OPEN,
            ltout => \N_1045_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_i_m2_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__15142\,
            in1 => \N__13004\,
            in2 => \N__12998\,
            in3 => \N__14087\,
            lcout => \N_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16339\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12964\,
            in2 => \N__12995\,
            in3 => \N__12986\,
            lcout => if_generate_plus_mult1_un68_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15413\,
            in2 => \N__12983\,
            in3 => \N__12968\,
            lcout => if_generate_plus_mult1_un68_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16003\,
            in1 => \N__12965\,
            in2 => \N__12956\,
            in3 => \N__12944\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_s_5_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12941\,
            in2 => \_gnd_net_\,
            in3 => \N__12932\,
            lcout => un5_rowlto2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_3_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001010"
        )
    port map (
            in0 => \N__12929\,
            in1 => \N__12923\,
            in2 => \N__12917\,
            in3 => \N__13076\,
            lcout => OPEN,
            ltout => \Pixel_1_r_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13193\,
            in2 => \N__13187\,
            in3 => \N__13184\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \m6_1_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000111100"
        )
    port map (
            in0 => \N__15414\,
            in1 => \N__15686\,
            in2 => \N__15873\,
            in3 => \N__16015\,
            lcout => \m6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI1M3Q1V2_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011000"
        )
    port map (
            in0 => \N__13064\,
            in1 => \N__13205\,
            in2 => \N__13325\,
            in3 => \N__14504\,
            lcout => OPEN,
            ltout => \beamX_RNI1M3Q1V2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIB75H7E_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13091\,
            in2 => \N__13079\,
            in3 => \N__13259\,
            lcout => \N_1039_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIAQ1S27_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__14533\,
            in1 => \N__14412\,
            in2 => \_gnd_net_\,
            in3 => \N__14578\,
            lcout => font_un3_pixel_29,
            ltout => \font_un3_pixel_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI440R9C_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101100110"
        )
    port map (
            in0 => \N__14579\,
            in1 => \N__14534\,
            in2 => \N__13070\,
            in3 => \N__14501\,
            lcout => OPEN,
            ltout => \G_7_0_m4_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNII9SNAB_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111010"
        )
    port map (
            in0 => \N__14502\,
            in1 => \N__14738\,
            in2 => \N__13067\,
            in3 => \N__14678\,
            lcout => \G_7_0_m4_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7OTDJ61_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__13058\,
            in1 => \_gnd_net_\,
            in2 => \N__15209\,
            in3 => \N__13375\,
            lcout => OPEN,
            ltout => \beamY_RNI7OTDJ61Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__font_un126_pixel_6_am_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__14535\,
            in1 => \N__14580\,
            in2 => \N__13049\,
            in3 => \N__13274\,
            lcout => OPEN,
            ltout => \font_un126_pixel_6_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIQ6MATS2_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14503\,
            in2 => \N__13268\,
            in3 => \N__13265\,
            lcout => \beamX_RNIQ6MATS2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII25UDD3_1_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__13249\,
            in1 => \N__15127\,
            in2 => \_gnd_net_\,
            in3 => \N__14381\,
            lcout => \beamY_RNII25UDD3_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m36_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__15841\,
            in1 => \N__16054\,
            in2 => \_gnd_net_\,
            in3 => \N__15673\,
            lcout => OPEN,
            ltout => \N_37_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI05CI5A3_1_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15128\,
            in2 => \N__13226\,
            in3 => \N__15176\,
            lcout => OPEN,
            ltout => \beamY_RNI05CI5A3_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJFRDMU2_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__13377\,
            in1 => \N__14654\,
            in2 => \N__13223\,
            in3 => \N__14937\,
            lcout => OPEN,
            ltout => \un116_pixel_7_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFHEQCT1_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__13220\,
            in1 => \N__13214\,
            in2 => \N__13208\,
            in3 => \N__13378\,
            lcout => \beamY_RNIFHEQCT1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIA4V0NM1_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000010"
        )
    port map (
            in0 => \N__15842\,
            in1 => \N__13280\,
            in2 => \N__15161\,
            in3 => \N__15674\,
            lcout => OPEN,
            ltout => \beamY_RNIA4V0NM1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUJBUM5_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__13286\,
            in1 => \N__14930\,
            in2 => \N__13196\,
            in3 => \N__13376\,
            lcout => OPEN,
            ltout => \un116_pixel_7_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBHJ7AM_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__14669\,
            in1 => \N__13400\,
            in2 => \N__13391\,
            in3 => \N__13381\,
            lcout => \beamY_RNIBHJ7AMZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16583\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13304\,
            in2 => \N__13316\,
            in3 => \N__15582\,
            lcout => \G_340\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13478\,
            in2 => \N__15657\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13298\,
            in2 => \N__13460\,
            in3 => \N__15583\,
            lcout => \G_341\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_s_5_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13448\,
            in2 => \_gnd_net_\,
            in3 => \N__13292\,
            lcout => un5_rowlto0,
            ltout => \un5_rowlto0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m39_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000100000"
        )
    port map (
            in0 => \N__15632\,
            in1 => \N__16035\,
            in2 => \N__13289\,
            in3 => \N__15475\,
            lcout => \un114_pixel_0_1__N_6_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJ720T72_0_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000110110010"
        )
    port map (
            in0 => \N__16037\,
            in1 => \N__13427\,
            in2 => \N__15163\,
            in3 => \N__15848\,
            lcout => \beamY_RNIJ720T72Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHD4CEK_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__15137\,
            in1 => \N__16036\,
            in2 => \_gnd_net_\,
            in3 => \N__15476\,
            lcout => un116_pixel_5_ns_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16454\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16094\,
            in2 => \N__13490\,
            in3 => \N__13472\,
            lcout => if_generate_plus_mult1_un75_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13469\,
            in2 => \N__16087\,
            in3 => \N__13451\,
            lcout => if_generate_plus_mult1_un75_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15587\,
            in1 => \N__13406\,
            in2 => \N__13421\,
            in3 => \N__13442\,
            lcout => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_s_5_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13439\,
            in2 => \_gnd_net_\,
            in3 => \N__13430\,
            lcout => un5_rowlto1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m2_0_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15588\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15467\,
            lcout => \N_321\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6CDEHM3_0_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001111111"
        )
    port map (
            in0 => \N__15468\,
            in1 => \N__15133\,
            in2 => \N__16088\,
            in3 => \N__15589\,
            lcout => un116_pixel_2_ns_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__13420\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16071\,
            lcout => if_generate_plus_mult1_un75_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14221\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIH_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13700\,
            in2 => \_gnd_net_\,
            in3 => \N__13760\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNIBVIHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13958\,
            in2 => \_gnd_net_\,
            in3 => \N__13542\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14222\,
            in2 => \_gnd_net_\,
            in3 => \N__13727\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRB_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14226\,
            in2 => \N__14265\,
            in3 => \N__13715\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI3HRBZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13706\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13703\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__SUM5_3_a3_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13682\,
            in2 => \_gnd_net_\,
            in3 => \N__13615\,
            lcout => \N_520\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13828\,
            in2 => \N__13508\,
            in3 => \N__13493\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13982\,
            in2 => \N__13816\,
            in3 => \N__13976\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI6FGK1_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13789\,
            in1 => \N__13829\,
            in2 => \N__13973\,
            in3 => \N__13964\,
            lcout => charx_if_generate_plus_mult1_un40_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13957\,
            in1 => \N__13841\,
            in2 => \N__13817\,
            in3 => \N__13835\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0\,
            ltout => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99QZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIK99Q_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13832\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13827\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14346\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONU_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13802\,
            in2 => \N__14074\,
            in3 => \N__13793\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNISONUZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRG1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13790\,
            in2 => \N__13778\,
            in3 => \N__13769\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIUPRGZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNI5LOD3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14012\,
            in1 => \N__13766\,
            in2 => \N__14075\,
            in3 => \N__14060\,
            lcout => charx_if_generate_plus_mult1_un47_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14057\,
            in2 => \_gnd_net_\,
            in3 => \N__14051\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTMZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15287\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URT1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14288\,
            in2 => \N__13996\,
            in3 => \N__14048\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI1URTZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQ2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14011\,
            in2 => \N__14045\,
            in3 => \N__14036\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNI3LHQZ0Z2\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI0GDV6_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16243\,
            in1 => \N__14033\,
            in2 => \N__13997\,
            in3 => \N__14027\,
            lcout => charx_if_generate_plus_mult1_un54_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14024\,
            in2 => \_gnd_net_\,
            in3 => \N__14018\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3\,
            ltout => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMIZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIQNMI3_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14015\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIKTTM1_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14010\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14351\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16466\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADB3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16664\,
            in3 => \N__14282\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNI1VADBZ0Z3\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14270\,
            in2 => \N__16652\,
            in3 => \N__14096\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16621\,
            in3 => \N__14093\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14090\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__g0_10_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000110011"
        )
    port map (
            in0 => \N__14536\,
            in1 => \N__14414\,
            in2 => \_gnd_net_\,
            in3 => \N__14581\,
            lcout => \un114_pixel_6_1_5__g2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14531\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TR1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14617\,
            in2 => \N__16598\,
            in3 => \N__14078\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI5Q8TRZ0Z1\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPB3_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14636\,
            in2 => \N__14599\,
            in3 => \N__14630\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIBLGPBZ0Z3\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14618\,
            in2 => \N__14627\,
            in3 => \N__14616\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPB3_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14606\,
            in1 => \N__16622\,
            in2 => \N__14600\,
            in3 => \N__14585\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3\,
            ltout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNIFTKPBZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__font_un126_pixel_m_1_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011111101101"
        )
    port map (
            in0 => \N__14532\,
            in1 => \N__14558\,
            in2 => \N__14552\,
            in3 => \N__14393\,
            lcout => \un114_pixel_6_1_5__font_un126_pixel_m_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIM245R1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16577\,
            in2 => \_gnd_net_\,
            in3 => \N__16499\,
            lcout => charx_if_generate_plus_mult1_un1_sum_axb1,
            ltout => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__font_un126_pixel_m_1_1_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011001010110"
        )
    port map (
            in0 => \N__14498\,
            in1 => \N__14413\,
            in2 => \N__14396\,
            in3 => \_gnd_net_\,
            lcout => \un114_pixel_6_1_5__font_un126_pixel_m_1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_4_0_15__m15_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100001100000"
        )
    port map (
            in0 => \N__15680\,
            in1 => \N__16011\,
            in2 => \N__15874\,
            in3 => \N__15495\,
            lcout => OPEN,
            ltout => \m15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII25UDD3_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__15146\,
            in1 => \_gnd_net_\,
            in2 => \N__14387\,
            in3 => \N__14384\,
            lcout => \beamY_RNII25UDD3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI4NRC8D1_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011010100"
        )
    port map (
            in0 => \N__16012\,
            in1 => \N__14663\,
            in2 => \N__15165\,
            in3 => \N__14724\,
            lcout => OPEN,
            ltout => \beamY_RNI4NRC8D1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNID79CMQ_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14925\,
            in2 => \N__14687\,
            in3 => \N__14684\,
            lcout => \N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBKJ0H51_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101000011"
        )
    port map (
            in0 => \N__15496\,
            in1 => \N__15868\,
            in2 => \N__15164\,
            in3 => \N__15681\,
            lcout => OPEN,
            ltout => \un116_pixel_2_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIH01F2S_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__14725\,
            in1 => \N__15153\,
            in2 => \N__14672\,
            in3 => \N__16013\,
            lcout => \beamY_RNIH01F2SZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_2_ns_1_5_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110011"
        )
    port map (
            in0 => \N__15492\,
            in1 => \N__15794\,
            in2 => \N__16085\,
            in3 => \N__15678\,
            lcout => \un116_pixel_2_ns_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__un114_pixel_3_0_3_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110111101101"
        )
    port map (
            in0 => \N__15679\,
            in1 => \N__16066\,
            in2 => \N__15852\,
            in3 => \N__15494\,
            lcout => OPEN,
            ltout => \N_276_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII25UDD3_3_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15109\,
            in2 => \N__14657\,
            in3 => \N__14645\,
            lcout => \beamY_RNII25UDD3_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m7_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100100100001"
        )
    port map (
            in0 => \N__15677\,
            in1 => \N__16061\,
            in2 => \N__15851\,
            in3 => \N__15491\,
            lcout => m7,
            ltout => \m7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNII25UDD3_2_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15108\,
            in2 => \N__14639\,
            in3 => \N__15193\,
            lcout => un116_pixel_3_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15493\,
            lcout => \N_302_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITQPUS72_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010010101"
        )
    port map (
            in0 => \N__16065\,
            in1 => \N__15182\,
            in2 => \N__15160\,
            in3 => \N__15793\,
            lcout => OPEN,
            ltout => \beamY_RNITQPUS72Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6B7UAL1_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__14924\,
            in1 => \_gnd_net_\,
            in2 => \N__15218\,
            in3 => \N__15215\,
            lcout => \beamY_RNI6B7UAL1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m31_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000000011"
        )
    port map (
            in0 => \N__15497\,
            in1 => \N__15624\,
            in2 => \N__15849\,
            in3 => \N__16056\,
            lcout => m31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_4_1_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101111"
        )
    port map (
            in0 => \N__16057\,
            in1 => \_gnd_net_\,
            in2 => \N__15675\,
            in3 => \N__15498\,
            lcout => \un116_pixel_4_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_6_1_5__m38_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__15500\,
            in1 => \N__15631\,
            in2 => \N__15850\,
            in3 => \N__16060\,
            lcout => m38,
            ltout => \m38_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPG8ISM3_1_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100011001"
        )
    port map (
            in0 => \N__14923\,
            in1 => \N__15138\,
            in2 => \N__14942\,
            in3 => \N__15789\,
            lcout => OPEN,
            ltout => \un116_pixel_6_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICKDGA43_1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__14938\,
            in1 => \N__14693\,
            in2 => \N__14741\,
            in3 => \N__15347\,
            lcout => \N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_2_bm_1_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__16058\,
            in1 => \N__14722\,
            in2 => \_gnd_net_\,
            in3 => \N__15788\,
            lcout => \un116_pixel_2_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_rowlto2_sbtinv_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16055\,
            lcout => un5_rowlto2_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_2_am_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010010110100"
        )
    port map (
            in0 => \N__16059\,
            in1 => \N__15787\,
            in2 => \N__15676\,
            in3 => \N__15499\,
            lcout => \un116_pixel_2_amZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16136\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQV3_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15239\,
            in2 => \N__15341\,
            in3 => \N__15326\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNI3UQVZ0Z3\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLR5_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15323\,
            in2 => \N__16253\,
            in3 => \N__15311\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNICTLRZ0Z5\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNI57HTG_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16216\,
            in1 => \N__16267\,
            in2 => \N__16229\,
            in3 => \N__15308\,
            lcout => charx_if_generate_plus_mult1_un61_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15305\,
            in2 => \_gnd_net_\,
            in3 => \N__15293\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7\,
            ltout => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIAZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIJRIA7_0_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15290\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8D6_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16268\,
            in2 => \_gnd_net_\,
            in3 => \N__16249\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNITC8DZ0Z6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16326\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TD7_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16100\,
            in2 => \N__16186\,
            in3 => \N__16220\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNIO7TDZ0Z7\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBB_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16217\,
            in2 => \N__16205\,
            in3 => \N__16196\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI5AOBBZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNI57I6U_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16399\,
            in1 => \N__16193\,
            in2 => \N__16187\,
            in3 => \N__16172\,
            lcout => charx_if_generate_plus_mult1_un68_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16169\,
            in2 => \_gnd_net_\,
            in3 => \N__16163\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0\,
            ltout => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUGZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNIMRTUG_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16160\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16155\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16447\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4H_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16295\,
            in2 => \N__16369\,
            in3 => \N__16403\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNI0PN4HZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGO_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16400\,
            in2 => \N__16388\,
            in3 => \N__16379\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNI48MGOZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNIFS1PQ1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16708\,
            in1 => \N__16376\,
            in2 => \N__16370\,
            in3 => \N__16355\,
            lcout => charx_if_generate_plus_mult1_un75_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAU_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16352\,
            in2 => \_gnd_net_\,
            in3 => \N__16346\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNITFFAUZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_0_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16327\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16562\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630C_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16289\,
            in2 => \N__16690\,
            in3 => \N__16280\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNI630CZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PF1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16277\,
            in2 => \N__16709\,
            in3 => \N__16271\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIHM9PFZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16715\,
            in2 => \N__16691\,
            in3 => \N__16704\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63R1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16676\,
            in3 => \N__16667\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNI5E63RZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000001111"
        )
    port map (
            in0 => \N__16579\,
            in1 => \N__16514\,
            in2 => \N__16639\,
            in3 => \N__16486\,
            lcout => charx_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_0_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000101111"
        )
    port map (
            in0 => \N__16515\,
            in1 => \N__16581\,
            in2 => \N__16495\,
            in3 => \N__16635\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNIDSDAB3_1_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111110000"
        )
    port map (
            in0 => \N__16580\,
            in1 => \N__16516\,
            in2 => \N__16640\,
            in3 => \N__16490\,
            lcout => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIS54HR1_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110100101"
        )
    port map (
            in0 => \N__16491\,
            in1 => \_gnd_net_\,
            in2 => \N__16520\,
            in3 => \N__16582\,
            lcout => charx_i_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__16578\,
            in1 => \N__16513\,
            in2 => \_gnd_net_\,
            in3 => \N__16485\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
