-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 17 2015 17:51:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSyncDebug : out std_logic;
    PixelDebug : out std_logic;
    HSyncDebug : out std_logic;
    Clock12MHz : in std_logic;
    VSync : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4347\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4263\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4002\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3957\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3867\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3753\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3504\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3495\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3489\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3317\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3287\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3249\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3141\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3090\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2916\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2766\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2757\ : std_logic;
signal \N__2754\ : std_logic;
signal \N__2751\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2691\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2672\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2670\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2666\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2648\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2645\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2552\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2486\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2459\ : std_logic;
signal \N__2456\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2432\ : std_logic;
signal \N__2429\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2414\ : std_logic;
signal \N__2411\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2399\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2378\ : std_logic;
signal \N__2375\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2349\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2346\ : std_logic;
signal \N__2343\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2288\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2252\ : std_logic;
signal \N__2249\ : std_logic;
signal \N__2246\ : std_logic;
signal \N__2243\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \VCCG0\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \Clock12MHz_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_7_1_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3UZ0\ : std_logic;
signal \bfn_7_2_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1FZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum_i\ : std_logic;
signal \un5_beamx_0_a2_3_cascade_\ : std_logic;
signal \un5_beamx_0_a2_5_cascade_\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal un5_beamx : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_i_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPFZ0Z3\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_axb_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum_i\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un47_sum\ : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un40_sum\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_8_4_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal \Pixel_0_sqmuxa_i_2_1_cascade_\ : std_logic;
signal \un1_beamylto9_0_a2_1_cascade_\ : std_logic;
signal \VSync_c\ : std_logic;
signal \N_84_cascade_\ : std_logic;
signal \N_132\ : std_logic;
signal \Pixel_0_sqmuxa_i_2\ : std_logic;
signal \N_101_cascade_\ : std_logic;
signal \Pixel_0_sqmuxa_i_1\ : std_logic;
signal un1_beamylto9_0_a2_1 : std_logic;
signal \Pixel_0_sqmuxa_i_4_cascade_\ : std_logic;
signal \N_99\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0_cascade_\ : std_logic;
signal \N_98\ : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal un5_visibley_cry_0 : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal un5_visibley_cry_1 : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal un5_visibley_cry_2 : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal un5_visibley_cry_3 : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal un5_visibley_cry_4 : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal un5_visibley_cry_5 : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal un5_visibley_cry_6 : std_logic;
signal un5_visibley_cry_7 : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal un5_visibley_cry_8 : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_i_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_axb_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un54_sum_i\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FEZ0Z21\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_i_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQEZ0Z1\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_axb_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un61_sum_i\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_i\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BKZ0Z1\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNKZ0Z2\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un68_sum_i_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_6\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_axb_8\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6_cascade_\ : std_logic;
signal \Pixel_1_RNOZ0Z_7\ : std_logic;
signal un5_visiblex_i : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0\ : std_logic;
signal \un5_visiblex_i_cascade_\ : std_logic;
signal \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6\ : std_logic;
signal un3_beamx_i_i_a2_4 : std_logic;
signal \un3_beamx_i_i_a2_5_cascade_\ : std_logic;
signal \beamX_RNI5457Z0Z_1\ : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal \N_97\ : std_logic;
signal \N_87\ : std_logic;
signal \N_130_cascade_\ : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal \HSync_c\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94_cascade_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVFZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GIZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6IIZ0Z1\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1_cascade_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum : std_logic;
signal un1_visibley_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PPZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULVZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_axb_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un26_sum : std_logic;
signal \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum : std_logic;
signal un1_visibley_if_generate_plus_mult1_un33_sum_i_0 : std_logic;
signal \un5_visibley_cry_0_c_RNIJVSBZ0\ : std_logic;
signal \N_8_cascade_\ : std_logic;
signal \Pixel_0_sqmuxa_i_5\ : std_logic;
signal \N_94\ : std_logic;
signal \N_49_cascade_\ : std_logic;
signal \N_59\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \Pixel_1_RNOZ0Z_6\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32\ : std_logic;
signal \G_7_0_a4_0_0\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32_cascade_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1\ : std_logic;
signal \N_11\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJIZ0Z2\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6PZ0Z3\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QORZ0Z3\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un47_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8_cascade_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPHZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85QZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPUZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum : std_logic;
signal \bfn_12_5_0_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQNZ0Z8\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TMZ0Z4\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCDZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICAZ0Z117\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMFZ0\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIILZ0Z78\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un54_sum_i_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0\ : std_logic;
signal \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0_cascade_\ : std_logic;
signal un1_visibley_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \PixelDebug_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \VSyncDebug_wire\ : std_logic;
signal \Clock12MHz_wire\ : std_logic;
signal \HSyncDebug_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    PixelDebug <= \PixelDebug_wire\;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    Pixel <= \Pixel_wire\;
    VSyncDebug <= \VSyncDebug_wire\;
    \Clock12MHz_wire\ <= Clock12MHz;
    HSyncDebug <= \HSyncDebug_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__2234\,
            RESETB => \N__4061\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \PixelDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4782\,
            DIN => \N__4781\,
            DOUT => \N__4780\,
            PACKAGEPIN => \PixelDebug_wire\
        );

    \PixelDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4782\,
            PADOUT => \N__4781\,
            PADIN => \N__4780\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4217\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4773\,
            DIN => \N__4772\,
            DOUT => \N__4771\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4773\,
            PADOUT => \N__4772\,
            PADIN => \N__4771\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2608\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4764\,
            DIN => \N__4763\,
            DOUT => \N__4762\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4764\,
            PADOUT => \N__4763\,
            PADIN => \N__4762\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4755\,
            DIN => \N__4754\,
            DOUT => \N__4753\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4755\,
            PADOUT => \N__4754\,
            PADIN => \N__4753\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4213\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4746\,
            DIN => \N__4745\,
            DOUT => \N__4744\,
            PACKAGEPIN => \VSyncDebug_wire\
        );

    \VSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4746\,
            PADOUT => \N__4745\,
            PADIN => \N__4744\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2618\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Clock12MHz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4737\,
            DIN => \N__4736\,
            DOUT => \N__4735\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4737\,
            PADOUT => \N__4736\,
            PADIN => \N__4735\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \Clock12MHz_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSyncDebug_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4728\,
            DIN => \N__4727\,
            DOUT => \N__4726\,
            PACKAGEPIN => \HSyncDebug_wire\
        );

    \HSyncDebug_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4728\,
            PADOUT => \N__4727\,
            PADIN => \N__4726\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3662\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1025\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4705\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4702\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__1021\ : Span4Mux_v
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__1020\ : Span4Mux_s3_h
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__4693\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__4690\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__4685\,
            I => \N__4682\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4679\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4679\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__1014\ : InMux
    port map (
            O => \N__4676\,
            I => \N__4673\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__4673\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQNZ0Z8\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4670\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__1011\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4664\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TMZ0Z4\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__4661\,
            I => \N__4658\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__4655\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCDZ0\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4652\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__4649\,
            I => \N__4645\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4636\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4636\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4636\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4633\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4636\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4633\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__997\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__4622\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICAZ0Z117\
        );

    \I__995\ : InMux
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4616\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMFZ0\
        );

    \I__993\ : InMux
    port map (
            O => \N__4613\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__992\ : InMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4607\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIILZ0Z78\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__989\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4598\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_i_7
        );

    \I__987\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4592\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__985\ : InMux
    port map (
            O => \N__4589\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__984\ : InMux
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4583\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__982\ : InMux
    port map (
            O => \N__4580\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__4577\,
            I => \N__4573\
        );

    \I__980\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4564\
        );

    \I__979\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4564\
        );

    \I__978\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4564\
        );

    \I__977\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4561\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4564\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4561\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__4556\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0_cascade_\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__972\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4547\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__4544\,
            I => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8_cascade_\
        );

    \I__969\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4535\
        );

    \I__968\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4535\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__966\ : Span4Mux_s3_h
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__4529\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum
        );

    \I__964\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4522\
        );

    \I__963\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4519\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__4522\,
            I => \N__4514\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4519\,
            I => \N__4514\
        );

    \I__960\ : Span4Mux_s3_h
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__959\ : Odrv4
    port map (
            O => \N__4511\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__957\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4502\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__4502\,
            I => \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPHZ0\
        );

    \I__955\ : InMux
    port map (
            O => \N__4499\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__954\ : InMux
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4493\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85QZ0\
        );

    \I__952\ : InMux
    port map (
            O => \N__4490\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__951\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4484\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4484\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPUZ0\
        );

    \I__949\ : InMux
    port map (
            O => \N__4481\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__947\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4472\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__945\ : InMux
    port map (
            O => \N__4469\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__944\ : InMux
    port map (
            O => \N__4466\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__4463\,
            I => \N__4458\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__4462\,
            I => \N__4454\
        );

    \I__941\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4450\
        );

    \I__940\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4441\
        );

    \I__939\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4441\
        );

    \I__938\ : InMux
    port map (
            O => \N__4454\,
            I => \N__4441\
        );

    \I__937\ : InMux
    port map (
            O => \N__4453\,
            I => \N__4441\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4450\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4441\,
            I => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__4436\,
            I => \N__4433\
        );

    \I__933\ : InMux
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4430\,
            I => un1_visibley_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__931\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__929\ : Odrv12
    port map (
            O => \N__4421\,
            I => \G_7_0_a4_0_0\
        );

    \I__928\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4414\
        );

    \I__927\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4411\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4414\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4411\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__4406\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32_cascade_\
        );

    \I__923\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4399\
        );

    \I__922\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4396\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4399\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4396\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1\
        );

    \I__919\ : InMux
    port map (
            O => \N__4391\,
            I => \N__4388\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__4388\,
            I => \N_11\
        );

    \I__917\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4382\,
            I => un1_visibley_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__914\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__4370\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__911\ : InMux
    port map (
            O => \N__4367\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__910\ : InMux
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__4358\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJIZ0Z2\
        );

    \I__907\ : InMux
    port map (
            O => \N__4355\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__4352\,
            I => \N__4348\
        );

    \I__905\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4340\
        );

    \I__904\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4340\
        );

    \I__903\ : InMux
    port map (
            O => \N__4347\,
            I => \N__4340\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4340\,
            I => \N__4336\
        );

    \I__901\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4333\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__4336\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__4333\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__897\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__4319\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6PZ0Z3\
        );

    \I__894\ : InMux
    port map (
            O => \N__4316\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__893\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__4307\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QORZ0Z3\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__889\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__4295\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_i_7
        );

    \I__886\ : InMux
    port map (
            O => \N__4292\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__885\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__4283\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__882\ : InMux
    port map (
            O => \N__4280\,
            I => un1_visibley_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__881\ : InMux
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4274\,
            I => \N__4269\
        );

    \I__879\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4266\
        );

    \I__878\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4263\
        );

    \I__877\ : Span4Mux_s3_h
    port map (
            O => \N__4269\,
            I => \N__4258\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4266\,
            I => \N__4258\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4263\,
            I => \un5_visibley_cry_0_c_RNIJVSBZ0\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__4258\,
            I => \un5_visibley_cry_0_c_RNIJVSBZ0\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__4253\,
            I => \N_8_cascade_\
        );

    \I__872\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4247\,
            I => \N__4244\
        );

    \I__870\ : Span4Mux_s3_h
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__4241\,
            I => \Pixel_0_sqmuxa_i_5\
        );

    \I__868\ : InMux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__4232\,
            I => \N_94\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__4229\,
            I => \N_49_cascade_\
        );

    \I__864\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__4220\,
            I => \N_59\
        );

    \I__861\ : IoInMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4214\,
            I => \N__4210\
        );

    \I__859\ : IoInMux
    port map (
            O => \N__4213\,
            I => \N__4207\
        );

    \I__858\ : Span4Mux_s2_v
    port map (
            O => \N__4210\,
            I => \N__4204\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4201\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4204\,
            I => \N__4198\
        );

    \I__855\ : IoSpan4Mux
    port map (
            O => \N__4201\,
            I => \N__4195\
        );

    \I__854\ : Span4Mux_v
    port map (
            O => \N__4198\,
            I => \N__4192\
        );

    \I__853\ : Span4Mux_s2_v
    port map (
            O => \N__4195\,
            I => \N__4189\
        );

    \I__852\ : Odrv4
    port map (
            O => \N__4192\,
            I => \Pixel_c\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__4189\,
            I => \Pixel_c\
        );

    \I__850\ : ClkMux
    port map (
            O => \N__4184\,
            I => \N__4160\
        );

    \I__849\ : ClkMux
    port map (
            O => \N__4183\,
            I => \N__4160\
        );

    \I__848\ : ClkMux
    port map (
            O => \N__4182\,
            I => \N__4160\
        );

    \I__847\ : ClkMux
    port map (
            O => \N__4181\,
            I => \N__4160\
        );

    \I__846\ : ClkMux
    port map (
            O => \N__4180\,
            I => \N__4160\
        );

    \I__845\ : ClkMux
    port map (
            O => \N__4179\,
            I => \N__4160\
        );

    \I__844\ : ClkMux
    port map (
            O => \N__4178\,
            I => \N__4160\
        );

    \I__843\ : ClkMux
    port map (
            O => \N__4177\,
            I => \N__4160\
        );

    \I__842\ : GlobalMux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__841\ : gio2CtrlBuf
    port map (
            O => \N__4157\,
            I => \PixelClock_g\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__839\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4146\
        );

    \I__838\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4143\
        );

    \I__837\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4140\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4146\,
            I => \N__4137\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4143\,
            I => \N__4132\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4132\
        );

    \I__833\ : Span4Mux_s3_h
    port map (
            O => \N__4137\,
            I => \N__4129\
        );

    \I__832\ : Span4Mux_s3_h
    port map (
            O => \N__4132\,
            I => \N__4126\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__4129\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum
        );

    \I__830\ : Odrv4
    port map (
            O => \N__4126\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum
        );

    \I__829\ : InMux
    port map (
            O => \N__4121\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__828\ : InMux
    port map (
            O => \N__4118\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__827\ : InMux
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4112\,
            I => \Pixel_1_RNOZ0Z_6\
        );

    \I__825\ : InMux
    port map (
            O => \N__4109\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__823\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4100\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4100\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\
        );

    \I__821\ : InMux
    port map (
            O => \N__4097\,
            I => un1_visibley_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__820\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4091\,
            I => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__817\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4082\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0\
        );

    \I__815\ : InMux
    port map (
            O => \N__4079\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__814\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4073\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0\
        );

    \I__812\ : InMux
    port map (
            O => \N__4070\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__811\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4064\,
            I => \un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PPZ0\
        );

    \I__809\ : IoInMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4058\,
            I => \N__4049\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4057\,
            I => \N__4046\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__4056\,
            I => \N__4043\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__4055\,
            I => \N__4040\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__4054\,
            I => \N__4037\
        );

    \I__803\ : InMux
    port map (
            O => \N__4053\,
            I => \N__4032\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__4052\,
            I => \N__4028\
        );

    \I__801\ : IoSpan4Mux
    port map (
            O => \N__4049\,
            I => \N__4025\
        );

    \I__800\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4020\
        );

    \I__799\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4020\
        );

    \I__798\ : InMux
    port map (
            O => \N__4040\,
            I => \N__4017\
        );

    \I__797\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4012\
        );

    \I__796\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4012\
        );

    \I__795\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4009\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4032\,
            I => \N__4006\
        );

    \I__793\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4003\
        );

    \I__792\ : InMux
    port map (
            O => \N__4028\,
            I => \N__3997\
        );

    \I__791\ : Span4Mux_s0_v
    port map (
            O => \N__4025\,
            I => \N__3994\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4020\,
            I => \N__3991\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4017\,
            I => \N__3986\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4012\,
            I => \N__3986\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__4009\,
            I => \N__3979\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__4006\,
            I => \N__3979\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4003\,
            I => \N__3979\
        );

    \I__784\ : InMux
    port map (
            O => \N__4002\,
            I => \N__3972\
        );

    \I__783\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3972\
        );

    \I__782\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3972\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__3997\,
            I => \N__3966\
        );

    \I__780\ : Span4Mux_v
    port map (
            O => \N__3994\,
            I => \N__3957\
        );

    \I__779\ : Span4Mux_v
    port map (
            O => \N__3991\,
            I => \N__3957\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__3986\,
            I => \N__3957\
        );

    \I__777\ : Span4Mux_v
    port map (
            O => \N__3979\,
            I => \N__3957\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3954\
        );

    \I__775\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3951\
        );

    \I__774\ : InMux
    port map (
            O => \N__3970\,
            I => \N__3946\
        );

    \I__773\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3946\
        );

    \I__772\ : Odrv12
    port map (
            O => \N__3966\,
            I => \CONSTANT_ONE_NET\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__3957\,
            I => \CONSTANT_ONE_NET\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__3954\,
            I => \CONSTANT_ONE_NET\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__3951\,
            I => \CONSTANT_ONE_NET\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3946\,
            I => \CONSTANT_ONE_NET\
        );

    \I__767\ : InMux
    port map (
            O => \N__3935\,
            I => \N__3932\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__3929\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULVZ0\
        );

    \I__764\ : InMux
    port map (
            O => \N__3926\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__3923\,
            I => \N__3919\
        );

    \I__762\ : InMux
    port map (
            O => \N__3922\,
            I => \N__3916\
        );

    \I__761\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3913\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__3916\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_axb_6
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3913\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_axb_6
        );

    \I__758\ : InMux
    port map (
            O => \N__3908\,
            I => \N__3905\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__3902\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\
        );

    \I__755\ : InMux
    port map (
            O => \N__3899\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__754\ : InMux
    port map (
            O => \N__3896\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_cry_6
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__3893\,
            I => \N__3890\
        );

    \I__752\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3887\,
            I => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO\
        );

    \I__750\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3877\
        );

    \I__749\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3877\
        );

    \I__748\ : InMux
    port map (
            O => \N__3882\,
            I => \N__3874\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3877\,
            I => \N__3867\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__3874\,
            I => \N__3867\
        );

    \I__745\ : InMux
    port map (
            O => \N__3873\,
            I => \N__3862\
        );

    \I__744\ : InMux
    port map (
            O => \N__3872\,
            I => \N__3862\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__3867\,
            I => un1_visibley_if_generate_plus_mult1_un26_sum
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3862\,
            I => un1_visibley_if_generate_plus_mult1_un26_sum
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__740\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3851\,
            I => \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\
        );

    \I__738\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3842\
        );

    \I__737\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3842\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3842\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum
        );

    \I__735\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3836\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__3836\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_i_0
        );

    \I__733\ : InMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__3830\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVFZ0Z1\
        );

    \I__731\ : InMux
    port map (
            O => \N__3827\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__3824\,
            I => \N__3821\
        );

    \I__729\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3818\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3818\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GIZ0Z1\
        );

    \I__727\ : InMux
    port map (
            O => \N__3815\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__726\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3809\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3809\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6IIZ0Z1\
        );

    \I__724\ : InMux
    port map (
            O => \N__3806\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__3803\,
            I => \N__3800\
        );

    \I__722\ : InMux
    port map (
            O => \N__3800\,
            I => \N__3797\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__3797\,
            I => un1_visibley_if_generate_plus_mult1_un33_sum_i_7
        );

    \I__720\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3791\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__3791\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_axb_7
        );

    \I__718\ : InMux
    port map (
            O => \N__3788\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__3785\,
            I => \N__3780\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__3784\,
            I => \N__3777\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__3783\,
            I => \N__3773\
        );

    \I__714\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3764\
        );

    \I__713\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3764\
        );

    \I__712\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3764\
        );

    \I__711\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3764\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__3764\,
            I => \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0\
        );

    \I__709\ : InMux
    port map (
            O => \N__3761\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__3758\,
            I => \N__3754\
        );

    \I__707\ : InMux
    port map (
            O => \N__3757\,
            I => \N__3745\
        );

    \I__706\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3745\
        );

    \I__705\ : InMux
    port map (
            O => \N__3753\,
            I => \N__3745\
        );

    \I__704\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3742\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3745\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__3742\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__3737\,
            I => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1_cascade_\
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__699\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3728\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__697\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3719\
        );

    \I__696\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3719\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__3719\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__693\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3710\,
            I => un1_visibley_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__691\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3700\
        );

    \I__690\ : InMux
    port map (
            O => \N__3706\,
            I => \N__3700\
        );

    \I__689\ : InMux
    port map (
            O => \N__3705\,
            I => \N__3697\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__3700\,
            I => \N_87\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__3697\,
            I => \N_87\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__3692\,
            I => \N_130_cascade_\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__3689\,
            I => \N__3683\
        );

    \I__684\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3680\
        );

    \I__683\ : InMux
    port map (
            O => \N__3687\,
            I => \N__3677\
        );

    \I__682\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3674\
        );

    \I__681\ : InMux
    port map (
            O => \N__3683\,
            I => \N__3671\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3680\,
            I => \beamXZ0Z_10\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3677\,
            I => \beamXZ0Z_10\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__3674\,
            I => \beamXZ0Z_10\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3671\,
            I => \beamXZ0Z_10\
        );

    \I__676\ : IoInMux
    port map (
            O => \N__3662\,
            I => \N__3659\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__674\ : IoSpan4Mux
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__673\ : Sp12to4
    port map (
            O => \N__3653\,
            I => \N__3649\
        );

    \I__672\ : IoInMux
    port map (
            O => \N__3652\,
            I => \N__3646\
        );

    \I__671\ : Span12Mux_v
    port map (
            O => \N__3649\,
            I => \N__3643\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3646\,
            I => \N__3640\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__3643\,
            I => \HSync_c\
        );

    \I__668\ : Odrv12
    port map (
            O => \N__3640\,
            I => \HSync_c\
        );

    \I__667\ : InMux
    port map (
            O => \N__3635\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__666\ : InMux
    port map (
            O => \N__3632\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__665\ : InMux
    port map (
            O => \N__3629\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__664\ : InMux
    port map (
            O => \N__3626\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__663\ : InMux
    port map (
            O => \N__3623\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__3620\,
            I => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94_cascade_\
        );

    \I__661\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3611\
        );

    \I__660\ : InMux
    port map (
            O => \N__3616\,
            I => \N__3611\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3611\,
            I => \N__3608\
        );

    \I__658\ : Odrv4
    port map (
            O => \N__3608\,
            I => un1_visibley_if_generate_plus_mult1_un47_sum
        );

    \I__657\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3602\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_axb_8\
        );

    \I__655\ : InMux
    port map (
            O => \N__3599\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__3596\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6_cascade_\
        );

    \I__653\ : InMux
    port map (
            O => \N__3593\,
            I => \N__3590\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3590\,
            I => \Pixel_1_RNOZ0Z_7\
        );

    \I__651\ : InMux
    port map (
            O => \N__3587\,
            I => \N__3578\
        );

    \I__650\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3578\
        );

    \I__649\ : InMux
    port map (
            O => \N__3585\,
            I => \N__3578\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3578\,
            I => un5_visiblex_i
        );

    \I__647\ : InMux
    port map (
            O => \N__3575\,
            I => \N__3569\
        );

    \I__646\ : InMux
    port map (
            O => \N__3574\,
            I => \N__3569\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3569\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__3566\,
            I => \un5_visiblex_i_cascade_\
        );

    \I__643\ : InMux
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3560\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6\
        );

    \I__641\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3554\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3554\,
            I => un3_beamx_i_i_a2_4
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__3551\,
            I => \un3_beamx_i_i_a2_5_cascade_\
        );

    \I__638\ : CEMux
    port map (
            O => \N__3548\,
            I => \N__3545\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3545\,
            I => \N__3540\
        );

    \I__636\ : CEMux
    port map (
            O => \N__3544\,
            I => \N__3537\
        );

    \I__635\ : CEMux
    port map (
            O => \N__3543\,
            I => \N__3533\
        );

    \I__634\ : Span4Mux_v
    port map (
            O => \N__3540\,
            I => \N__3528\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3537\,
            I => \N__3528\
        );

    \I__632\ : InMux
    port map (
            O => \N__3536\,
            I => \N__3525\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3533\,
            I => \N__3520\
        );

    \I__630\ : Span4Mux_h
    port map (
            O => \N__3528\,
            I => \N__3517\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3525\,
            I => \N__3514\
        );

    \I__628\ : InMux
    port map (
            O => \N__3524\,
            I => \N__3509\
        );

    \I__627\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3509\
        );

    \I__626\ : Span4Mux_v
    port map (
            O => \N__3520\,
            I => \N__3504\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__3517\,
            I => \N__3504\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__3514\,
            I => \beamX_RNI5457Z0Z_1\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3509\,
            I => \beamX_RNI5457Z0Z_1\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__3504\,
            I => \beamX_RNI5457Z0Z_1\
        );

    \I__621\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3490\
        );

    \I__620\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3486\
        );

    \I__619\ : InMux
    port map (
            O => \N__3495\,
            I => \N__3481\
        );

    \I__618\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3481\
        );

    \I__617\ : InMux
    port map (
            O => \N__3493\,
            I => \N__3478\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3490\,
            I => \N__3475\
        );

    \I__615\ : InMux
    port map (
            O => \N__3489\,
            I => \N__3472\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3486\,
            I => \beamXZ0Z_4\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3481\,
            I => \beamXZ0Z_4\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3478\,
            I => \beamXZ0Z_4\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__3475\,
            I => \beamXZ0Z_4\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__3472\,
            I => \beamXZ0Z_4\
        );

    \I__609\ : CascadeMux
    port map (
            O => \N__3461\,
            I => \N__3455\
        );

    \I__608\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3451\
        );

    \I__607\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3448\
        );

    \I__606\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3445\
        );

    \I__605\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3442\
        );

    \I__604\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3439\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3451\,
            I => \beamXZ0Z_6\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3448\,
            I => \beamXZ0Z_6\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3445\,
            I => \beamXZ0Z_6\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3442\,
            I => \beamXZ0Z_6\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3439\,
            I => \beamXZ0Z_6\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__3428\,
            I => \N__3424\
        );

    \I__597\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3418\
        );

    \I__596\ : InMux
    port map (
            O => \N__3424\,
            I => \N__3413\
        );

    \I__595\ : InMux
    port map (
            O => \N__3423\,
            I => \N__3413\
        );

    \I__594\ : InMux
    port map (
            O => \N__3422\,
            I => \N__3410\
        );

    \I__593\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3407\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__3418\,
            I => \beamXZ0Z_5\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__3413\,
            I => \beamXZ0Z_5\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3410\,
            I => \beamXZ0Z_5\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3407\,
            I => \beamXZ0Z_5\
        );

    \I__588\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3394\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__3397\,
            I => \N__3389\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3394\,
            I => \N__3386\
        );

    \I__585\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3383\
        );

    \I__584\ : InMux
    port map (
            O => \N__3392\,
            I => \N__3378\
        );

    \I__583\ : InMux
    port map (
            O => \N__3389\,
            I => \N__3378\
        );

    \I__582\ : Odrv4
    port map (
            O => \N__3386\,
            I => \N_97\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3383\,
            I => \N_97\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3378\,
            I => \N_97\
        );

    \I__579\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3367\
        );

    \I__578\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3364\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3367\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__3364\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__3359\,
            I => \N__3356\
        );

    \I__574\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3353\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3353\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FEZ0Z21\
        );

    \I__572\ : InMux
    port map (
            O => \N__3350\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\
        );

    \I__571\ : InMux
    port map (
            O => \N__3347\,
            I => \N__3341\
        );

    \I__570\ : InMux
    port map (
            O => \N__3346\,
            I => \N__3341\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3341\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_i_8\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__3338\,
            I => \N__3335\
        );

    \I__567\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3332\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3332\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQEZ0Z1\
        );

    \I__565\ : InMux
    port map (
            O => \N__3329\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\
        );

    \I__564\ : InMux
    port map (
            O => \N__3326\,
            I => \N__3323\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3323\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_axb_8\
        );

    \I__562\ : InMux
    port map (
            O => \N__3320\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7\
        );

    \I__561\ : InMux
    port map (
            O => \N__3317\,
            I => \N__3313\
        );

    \I__560\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3310\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3313\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3310\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__3305\,
            I => \N__3302\
        );

    \I__556\ : InMux
    port map (
            O => \N__3302\,
            I => \N__3299\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3299\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_i\
        );

    \I__554\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3290\
        );

    \I__553\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3290\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3290\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__3287\,
            I => \N__3284\
        );

    \I__550\ : InMux
    port map (
            O => \N__3284\,
            I => \N__3281\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3281\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_i\
        );

    \I__548\ : InMux
    port map (
            O => \N__3278\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\
        );

    \I__547\ : InMux
    port map (
            O => \N__3275\,
            I => \N__3272\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3272\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BKZ0Z1\
        );

    \I__545\ : InMux
    port map (
            O => \N__3269\,
            I => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3266\,
            I => \N__3263\
        );

    \I__543\ : InMux
    port map (
            O => \N__3263\,
            I => \N__3260\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__3260\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNKZ0Z2\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__3257\,
            I => \N__3253\
        );

    \I__540\ : InMux
    port map (
            O => \N__3256\,
            I => \N__3249\
        );

    \I__539\ : InMux
    port map (
            O => \N__3253\,
            I => \N__3244\
        );

    \I__538\ : InMux
    port map (
            O => \N__3252\,
            I => \N__3244\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__3249\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3244\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843\
        );

    \I__535\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3233\
        );

    \I__534\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3233\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3233\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_i_8\
        );

    \I__532\ : InMux
    port map (
            O => \N__3230\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\
        );

    \I__531\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3223\
        );

    \I__530\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3220\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3223\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3220\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__526\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3209\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3209\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0\
        );

    \I__524\ : InMux
    port map (
            O => \N__3206\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\
        );

    \I__523\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3197\
        );

    \I__522\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3197\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3197\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_i_8\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__3194\,
            I => \N__3191\
        );

    \I__519\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3188\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3188\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0\
        );

    \I__517\ : InMux
    port map (
            O => \N__3185\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\
        );

    \I__516\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3179\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3179\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_axb_8\
        );

    \I__514\ : InMux
    port map (
            O => \N__3176\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__3173\,
            I => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1_cascade_\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__3170\,
            I => \N__3166\
        );

    \I__511\ : InMux
    port map (
            O => \N__3169\,
            I => \N__3163\
        );

    \I__510\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3160\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3163\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3160\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__3155\,
            I => \N__3152\
        );

    \I__506\ : InMux
    port map (
            O => \N__3152\,
            I => \N__3149\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3149\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_i\
        );

    \I__504\ : InMux
    port map (
            O => \N__3146\,
            I => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\
        );

    \I__503\ : InMux
    port map (
            O => \N__3143\,
            I => \N__3134\
        );

    \I__502\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3134\
        );

    \I__501\ : InMux
    port map (
            O => \N__3141\,
            I => \N__3134\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3134\,
            I => \N__3128\
        );

    \I__499\ : InMux
    port map (
            O => \N__3133\,
            I => \N__3125\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__3132\,
            I => \N__3122\
        );

    \I__497\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3119\
        );

    \I__496\ : Span4Mux_h
    port map (
            O => \N__3128\,
            I => \N__3116\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3125\,
            I => \N__3113\
        );

    \I__494\ : InMux
    port map (
            O => \N__3122\,
            I => \N__3110\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3119\,
            I => \beamYZ0Z_2\
        );

    \I__492\ : Odrv4
    port map (
            O => \N__3116\,
            I => \beamYZ0Z_2\
        );

    \I__491\ : Odrv4
    port map (
            O => \N__3113\,
            I => \beamYZ0Z_2\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3110\,
            I => \beamYZ0Z_2\
        );

    \I__489\ : InMux
    port map (
            O => \N__3101\,
            I => un5_visibley_cry_1
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3098\,
            I => \N__3093\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__3097\,
            I => \N__3090\
        );

    \I__486\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3085\
        );

    \I__485\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3082\
        );

    \I__484\ : InMux
    port map (
            O => \N__3090\,
            I => \N__3079\
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__3089\,
            I => \N__3076\
        );

    \I__482\ : InMux
    port map (
            O => \N__3088\,
            I => \N__3073\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3085\,
            I => \N__3070\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3082\,
            I => \N__3065\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__3079\,
            I => \N__3065\
        );

    \I__478\ : InMux
    port map (
            O => \N__3076\,
            I => \N__3062\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3073\,
            I => \beamYZ0Z_3\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__3070\,
            I => \beamYZ0Z_3\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__3065\,
            I => \beamYZ0Z_3\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3062\,
            I => \beamYZ0Z_3\
        );

    \I__473\ : InMux
    port map (
            O => \N__3053\,
            I => un5_visibley_cry_2
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__3050\,
            I => \N__3046\
        );

    \I__471\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3041\
        );

    \I__470\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3038\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__3045\,
            I => \N__3034\
        );

    \I__468\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3031\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3041\,
            I => \N__3028\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3038\,
            I => \N__3025\
        );

    \I__465\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3022\
        );

    \I__464\ : InMux
    port map (
            O => \N__3034\,
            I => \N__3019\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__3031\,
            I => \beamYZ0Z_4\
        );

    \I__462\ : Odrv4
    port map (
            O => \N__3028\,
            I => \beamYZ0Z_4\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__3025\,
            I => \beamYZ0Z_4\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3022\,
            I => \beamYZ0Z_4\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3019\,
            I => \beamYZ0Z_4\
        );

    \I__458\ : InMux
    port map (
            O => \N__3008\,
            I => un5_visibley_cry_3
        );

    \I__457\ : InMux
    port map (
            O => \N__3005\,
            I => \N__2999\
        );

    \I__456\ : InMux
    port map (
            O => \N__3004\,
            I => \N__2996\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__3003\,
            I => \N__2992\
        );

    \I__454\ : InMux
    port map (
            O => \N__3002\,
            I => \N__2989\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2999\,
            I => \N__2986\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2996\,
            I => \N__2983\
        );

    \I__451\ : InMux
    port map (
            O => \N__2995\,
            I => \N__2980\
        );

    \I__450\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2977\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2989\,
            I => \beamYZ0Z_5\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__2986\,
            I => \beamYZ0Z_5\
        );

    \I__447\ : Odrv4
    port map (
            O => \N__2983\,
            I => \beamYZ0Z_5\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__2980\,
            I => \beamYZ0Z_5\
        );

    \I__445\ : LocalMux
    port map (
            O => \N__2977\,
            I => \beamYZ0Z_5\
        );

    \I__444\ : InMux
    port map (
            O => \N__2966\,
            I => un5_visibley_cry_4
        );

    \I__443\ : InMux
    port map (
            O => \N__2963\,
            I => \N__2958\
        );

    \I__442\ : InMux
    port map (
            O => \N__2962\,
            I => \N__2955\
        );

    \I__441\ : InMux
    port map (
            O => \N__2961\,
            I => \N__2950\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2958\,
            I => \N__2945\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2955\,
            I => \N__2945\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__2954\,
            I => \N__2942\
        );

    \I__437\ : InMux
    port map (
            O => \N__2953\,
            I => \N__2939\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__2950\,
            I => \N__2936\
        );

    \I__435\ : Span4Mux_h
    port map (
            O => \N__2945\,
            I => \N__2933\
        );

    \I__434\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2930\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2939\,
            I => \beamYZ0Z_6\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__2936\,
            I => \beamYZ0Z_6\
        );

    \I__431\ : Odrv4
    port map (
            O => \N__2933\,
            I => \beamYZ0Z_6\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2930\,
            I => \beamYZ0Z_6\
        );

    \I__429\ : InMux
    port map (
            O => \N__2921\,
            I => un5_visibley_cry_5
        );

    \I__428\ : InMux
    port map (
            O => \N__2918\,
            I => \N__2912\
        );

    \I__427\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2909\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__2916\,
            I => \N__2906\
        );

    \I__425\ : InMux
    port map (
            O => \N__2915\,
            I => \N__2903\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2912\,
            I => \N__2898\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2909\,
            I => \N__2898\
        );

    \I__422\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2895\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2903\,
            I => \beamYZ0Z_7\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__2898\,
            I => \beamYZ0Z_7\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2895\,
            I => \beamYZ0Z_7\
        );

    \I__418\ : InMux
    port map (
            O => \N__2888\,
            I => un5_visibley_cry_6
        );

    \I__417\ : InMux
    port map (
            O => \N__2885\,
            I => \N__2878\
        );

    \I__416\ : InMux
    port map (
            O => \N__2884\,
            I => \N__2873\
        );

    \I__415\ : InMux
    port map (
            O => \N__2883\,
            I => \N__2873\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__2882\,
            I => \N__2870\
        );

    \I__413\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2867\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2878\,
            I => \N__2862\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2873\,
            I => \N__2862\
        );

    \I__410\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2859\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__2867\,
            I => \beamYZ0Z_8\
        );

    \I__408\ : Odrv4
    port map (
            O => \N__2862\,
            I => \beamYZ0Z_8\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2859\,
            I => \beamYZ0Z_8\
        );

    \I__406\ : InMux
    port map (
            O => \N__2852\,
            I => \bfn_8_8_0_\
        );

    \I__405\ : InMux
    port map (
            O => \N__2849\,
            I => \N__2843\
        );

    \I__404\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2840\
        );

    \I__403\ : InMux
    port map (
            O => \N__2847\,
            I => \N__2837\
        );

    \I__402\ : InMux
    port map (
            O => \N__2846\,
            I => \N__2833\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2843\,
            I => \N__2828\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2840\,
            I => \N__2828\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2837\,
            I => \N__2825\
        );

    \I__398\ : InMux
    port map (
            O => \N__2836\,
            I => \N__2822\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2833\,
            I => \beamYZ0Z_9\
        );

    \I__396\ : Odrv4
    port map (
            O => \N__2828\,
            I => \beamYZ0Z_9\
        );

    \I__395\ : Odrv4
    port map (
            O => \N__2825\,
            I => \beamYZ0Z_9\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__2822\,
            I => \beamYZ0Z_9\
        );

    \I__393\ : InMux
    port map (
            O => \N__2813\,
            I => un5_visibley_cry_8
        );

    \I__392\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2807\,
            I => un1_beamylto9_0_a2_1
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__2804\,
            I => \Pixel_0_sqmuxa_i_4_cascade_\
        );

    \I__389\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2798\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__2798\,
            I => \N_99\
        );

    \I__387\ : InMux
    port map (
            O => \N__2795\,
            I => un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0
        );

    \I__386\ : InMux
    port map (
            O => \N__2792\,
            I => un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0
        );

    \I__385\ : InMux
    port map (
            O => \N__2789\,
            I => un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0
        );

    \I__384\ : CascadeMux
    port map (
            O => \N__2786\,
            I => \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0_cascade_\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__2783\,
            I => \N__2779\
        );

    \I__382\ : InMux
    port map (
            O => \N__2782\,
            I => \N__2774\
        );

    \I__381\ : InMux
    port map (
            O => \N__2779\,
            I => \N__2774\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2774\,
            I => \N_98\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__2771\,
            I => \N__2766\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__2770\,
            I => \N__2760\
        );

    \I__377\ : InMux
    port map (
            O => \N__2769\,
            I => \N__2757\
        );

    \I__376\ : InMux
    port map (
            O => \N__2766\,
            I => \N__2754\
        );

    \I__375\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2751\
        );

    \I__374\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2746\
        );

    \I__373\ : InMux
    port map (
            O => \N__2763\,
            I => \N__2746\
        );

    \I__372\ : InMux
    port map (
            O => \N__2760\,
            I => \N__2743\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__2757\,
            I => \beamYZ0Z_0\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2754\,
            I => \beamYZ0Z_0\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__2751\,
            I => \beamYZ0Z_0\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2746\,
            I => \beamYZ0Z_0\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2743\,
            I => \beamYZ0Z_0\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__2732\,
            I => \N__2724\
        );

    \I__365\ : InMux
    port map (
            O => \N__2731\,
            I => \N__2721\
        );

    \I__364\ : InMux
    port map (
            O => \N__2730\,
            I => \N__2718\
        );

    \I__363\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2713\
        );

    \I__362\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2713\
        );

    \I__361\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2710\
        );

    \I__360\ : InMux
    port map (
            O => \N__2724\,
            I => \N__2707\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2721\,
            I => \beamYZ0Z_1\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2718\,
            I => \beamYZ0Z_1\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2713\,
            I => \beamYZ0Z_1\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__2710\,
            I => \beamYZ0Z_1\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2707\,
            I => \beamYZ0Z_1\
        );

    \I__354\ : InMux
    port map (
            O => \N__2696\,
            I => un5_visibley_cry_0
        );

    \I__353\ : InMux
    port map (
            O => \N__2693\,
            I => \N__2687\
        );

    \I__352\ : InMux
    port map (
            O => \N__2692\,
            I => \N__2682\
        );

    \I__351\ : InMux
    port map (
            O => \N__2691\,
            I => \N__2682\
        );

    \I__350\ : InMux
    port map (
            O => \N__2690\,
            I => \N__2679\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2687\,
            I => \beamXZ0Z_7\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__2682\,
            I => \beamXZ0Z_7\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2679\,
            I => \beamXZ0Z_7\
        );

    \I__346\ : InMux
    port map (
            O => \N__2672\,
            I => \N__2666\
        );

    \I__345\ : InMux
    port map (
            O => \N__2671\,
            I => \N__2663\
        );

    \I__344\ : InMux
    port map (
            O => \N__2670\,
            I => \N__2660\
        );

    \I__343\ : InMux
    port map (
            O => \N__2669\,
            I => \N__2657\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2666\,
            I => \beamXZ0Z_8\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__2663\,
            I => \beamXZ0Z_8\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__2660\,
            I => \beamXZ0Z_8\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2657\,
            I => \beamXZ0Z_8\
        );

    \I__338\ : InMux
    port map (
            O => \N__2648\,
            I => \N__2641\
        );

    \I__337\ : InMux
    port map (
            O => \N__2647\,
            I => \N__2632\
        );

    \I__336\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2632\
        );

    \I__335\ : InMux
    port map (
            O => \N__2645\,
            I => \N__2632\
        );

    \I__334\ : InMux
    port map (
            O => \N__2644\,
            I => \N__2632\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2641\,
            I => \N__2629\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2632\,
            I => \beamXZ0Z_9\
        );

    \I__331\ : Odrv4
    port map (
            O => \N__2629\,
            I => \beamXZ0Z_9\
        );

    \I__330\ : CascadeMux
    port map (
            O => \N__2624\,
            I => \Pixel_0_sqmuxa_i_2_1_cascade_\
        );

    \I__329\ : CascadeMux
    port map (
            O => \N__2621\,
            I => \un1_beamylto9_0_a2_1_cascade_\
        );

    \I__328\ : IoInMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2615\,
            I => \N__2612\
        );

    \I__326\ : IoSpan4Mux
    port map (
            O => \N__2612\,
            I => \N__2609\
        );

    \I__325\ : Span4Mux_s1_v
    port map (
            O => \N__2609\,
            I => \N__2605\
        );

    \I__324\ : IoInMux
    port map (
            O => \N__2608\,
            I => \N__2602\
        );

    \I__323\ : Sp12to4
    port map (
            O => \N__2605\,
            I => \N__2599\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2602\,
            I => \N__2596\
        );

    \I__321\ : Odrv12
    port map (
            O => \N__2599\,
            I => \VSync_c\
        );

    \I__320\ : Odrv12
    port map (
            O => \N__2596\,
            I => \VSync_c\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__2591\,
            I => \N_84_cascade_\
        );

    \I__318\ : InMux
    port map (
            O => \N__2588\,
            I => \N__2584\
        );

    \I__317\ : InMux
    port map (
            O => \N__2587\,
            I => \N__2581\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__2584\,
            I => \N_132\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__2581\,
            I => \N_132\
        );

    \I__314\ : InMux
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__2573\,
            I => \Pixel_0_sqmuxa_i_2\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__2570\,
            I => \N_101_cascade_\
        );

    \I__311\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2564\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2564\,
            I => \Pixel_0_sqmuxa_i_1\
        );

    \I__309\ : InMux
    port map (
            O => \N__2561\,
            I => un8_beamx_cry_5
        );

    \I__308\ : InMux
    port map (
            O => \N__2558\,
            I => un8_beamx_cry_6
        );

    \I__307\ : InMux
    port map (
            O => \N__2555\,
            I => un8_beamx_cry_7
        );

    \I__306\ : InMux
    port map (
            O => \N__2552\,
            I => \bfn_8_4_0_\
        );

    \I__305\ : InMux
    port map (
            O => \N__2549\,
            I => un8_beamx_cry_9
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2546\,
            I => \N__2542\
        );

    \I__303\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2539\
        );

    \I__302\ : InMux
    port map (
            O => \N__2542\,
            I => \N__2536\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2539\,
            I => \beamXZ0Z_2\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2536\,
            I => \beamXZ0Z_2\
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__2531\,
            I => \N__2528\
        );

    \I__298\ : InMux
    port map (
            O => \N__2528\,
            I => \N__2525\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2525\,
            I => \N__2520\
        );

    \I__296\ : InMux
    port map (
            O => \N__2524\,
            I => \N__2515\
        );

    \I__295\ : InMux
    port map (
            O => \N__2523\,
            I => \N__2515\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__2520\,
            I => \beamXZ0Z_1\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2515\,
            I => \beamXZ0Z_1\
        );

    \I__292\ : InMux
    port map (
            O => \N__2510\,
            I => \N__2504\
        );

    \I__291\ : InMux
    port map (
            O => \N__2509\,
            I => \N__2497\
        );

    \I__290\ : InMux
    port map (
            O => \N__2508\,
            I => \N__2497\
        );

    \I__289\ : InMux
    port map (
            O => \N__2507\,
            I => \N__2497\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2504\,
            I => \beamXZ0Z_0\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2497\,
            I => \beamXZ0Z_0\
        );

    \I__286\ : InMux
    port map (
            O => \N__2492\,
            I => un5_visiblex_cry_5
        );

    \I__285\ : InMux
    port map (
            O => \N__2489\,
            I => un5_visiblex_cry_6
        );

    \I__284\ : InMux
    port map (
            O => \N__2486\,
            I => \N__2482\
        );

    \I__283\ : InMux
    port map (
            O => \N__2485\,
            I => \N__2479\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2482\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2479\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum\
        );

    \I__280\ : InMux
    port map (
            O => \N__2474\,
            I => un5_visiblex_cry_7
        );

    \I__279\ : InMux
    port map (
            O => \N__2471\,
            I => un5_visiblex_cry_8
        );

    \I__278\ : InMux
    port map (
            O => \N__2468\,
            I => \N__2462\
        );

    \I__277\ : InMux
    port map (
            O => \N__2467\,
            I => \N__2462\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2462\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum\
        );

    \I__275\ : InMux
    port map (
            O => \N__2459\,
            I => un8_beamx_cry_1
        );

    \I__274\ : InMux
    port map (
            O => \N__2456\,
            I => un8_beamx_cry_2
        );

    \I__273\ : InMux
    port map (
            O => \N__2453\,
            I => un8_beamx_cry_3
        );

    \I__272\ : InMux
    port map (
            O => \N__2450\,
            I => un8_beamx_cry_4
        );

    \I__271\ : InMux
    port map (
            O => \N__2447\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\
        );

    \I__270\ : InMux
    port map (
            O => \N__2444\,
            I => \N__2440\
        );

    \I__269\ : InMux
    port map (
            O => \N__2443\,
            I => \N__2437\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2440\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2437\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__2432\,
            I => \N__2429\
        );

    \I__265\ : InMux
    port map (
            O => \N__2429\,
            I => \N__2426\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2426\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365\
        );

    \I__263\ : InMux
    port map (
            O => \N__2423\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\
        );

    \I__262\ : InMux
    port map (
            O => \N__2420\,
            I => \N__2414\
        );

    \I__261\ : InMux
    port map (
            O => \N__2419\,
            I => \N__2414\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2414\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_i_8\
        );

    \I__259\ : CascadeMux
    port map (
            O => \N__2411\,
            I => \N__2408\
        );

    \I__258\ : InMux
    port map (
            O => \N__2408\,
            I => \N__2405\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2405\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPFZ0Z3\
        );

    \I__256\ : InMux
    port map (
            O => \N__2402\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\
        );

    \I__255\ : InMux
    port map (
            O => \N__2399\,
            I => \N__2396\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2396\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_axb_8\
        );

    \I__253\ : InMux
    port map (
            O => \N__2393\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7\
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__2390\,
            I => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0_cascade_\
        );

    \I__251\ : CascadeMux
    port map (
            O => \N__2387\,
            I => \N__2384\
        );

    \I__250\ : InMux
    port map (
            O => \N__2384\,
            I => \N__2381\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2381\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_i\
        );

    \I__248\ : InMux
    port map (
            O => \N__2378\,
            I => un5_visiblex_cry_4
        );

    \I__247\ : InMux
    port map (
            O => \N__2375\,
            I => un21_beamy_cry_1
        );

    \I__246\ : InMux
    port map (
            O => \N__2372\,
            I => un21_beamy_cry_2
        );

    \I__245\ : InMux
    port map (
            O => \N__2369\,
            I => un21_beamy_cry_3
        );

    \I__244\ : InMux
    port map (
            O => \N__2366\,
            I => un21_beamy_cry_4
        );

    \I__243\ : InMux
    port map (
            O => \N__2363\,
            I => un21_beamy_cry_5
        );

    \I__242\ : InMux
    port map (
            O => \N__2360\,
            I => un21_beamy_cry_6
        );

    \I__241\ : InMux
    port map (
            O => \N__2357\,
            I => un21_beamy_cry_7
        );

    \I__240\ : InMux
    port map (
            O => \N__2354\,
            I => \N__2350\
        );

    \I__239\ : InMux
    port map (
            O => \N__2353\,
            I => \N__2343\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2350\,
            I => \N__2340\
        );

    \I__237\ : InMux
    port map (
            O => \N__2349\,
            I => \N__2335\
        );

    \I__236\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2335\
        );

    \I__235\ : InMux
    port map (
            O => \N__2347\,
            I => \N__2330\
        );

    \I__234\ : InMux
    port map (
            O => \N__2346\,
            I => \N__2330\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2343\,
            I => \N__2327\
        );

    \I__232\ : Span4Mux_h
    port map (
            O => \N__2340\,
            I => \N__2322\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__2335\,
            I => \N__2322\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2330\,
            I => un5_beamx
        );

    \I__229\ : Odrv4
    port map (
            O => \N__2327\,
            I => un5_beamx
        );

    \I__228\ : Odrv4
    port map (
            O => \N__2322\,
            I => un5_beamx
        );

    \I__227\ : InMux
    port map (
            O => \N__2315\,
            I => \bfn_7_8_0_\
        );

    \I__226\ : CascadeMux
    port map (
            O => \N__2312\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\
        );

    \I__225\ : InMux
    port map (
            O => \N__2309\,
            I => \N__2306\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2306\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1FZ0\
        );

    \I__223\ : InMux
    port map (
            O => \N__2303\,
            I => \N__2300\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2300\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_i\
        );

    \I__221\ : CascadeMux
    port map (
            O => \N__2297\,
            I => \un5_beamx_0_a2_3_cascade_\
        );

    \I__220\ : CascadeMux
    port map (
            O => \N__2294\,
            I => \un5_beamx_0_a2_5_cascade_\
        );

    \I__219\ : InMux
    port map (
            O => \N__2291\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\
        );

    \I__218\ : InMux
    port map (
            O => \N__2288\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\
        );

    \I__217\ : InMux
    port map (
            O => \N__2285\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\
        );

    \I__216\ : InMux
    port map (
            O => \N__2282\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7\
        );

    \I__215\ : CascadeMux
    port map (
            O => \N__2279\,
            I => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_\
        );

    \I__214\ : CascadeMux
    port map (
            O => \N__2276\,
            I => \N__2273\
        );

    \I__213\ : InMux
    port map (
            O => \N__2273\,
            I => \N__2270\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__2270\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3UZ0\
        );

    \I__211\ : InMux
    port map (
            O => \N__2267\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5\
        );

    \I__210\ : InMux
    port map (
            O => \N__2264\,
            I => \N__2255\
        );

    \I__209\ : InMux
    port map (
            O => \N__2263\,
            I => \N__2255\
        );

    \I__208\ : InMux
    port map (
            O => \N__2262\,
            I => \N__2255\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__2255\,
            I => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__206\ : IoInMux
    port map (
            O => \N__2252\,
            I => \N__2249\
        );

    \I__205\ : LocalMux
    port map (
            O => \N__2249\,
            I => \N__2246\
        );

    \I__204\ : Span4Mux_s1_h
    port map (
            O => \N__2246\,
            I => \N__2243\
        );

    \I__203\ : Span4Mux_h
    port map (
            O => \N__2243\,
            I => \N__2240\
        );

    \I__202\ : Sp12to4
    port map (
            O => \N__2240\,
            I => \N__2237\
        );

    \I__201\ : Odrv12
    port map (
            O => \N__2237\,
            I => \Clock50MHz.PixelClock\
        );

    \I__200\ : IoInMux
    port map (
            O => \N__2234\,
            I => \N__2231\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__2231\,
            I => \N__2228\
        );

    \I__198\ : IoSpan4Mux
    port map (
            O => \N__2228\,
            I => \N__2225\
        );

    \I__197\ : Odrv4
    port map (
            O => \N__2225\,
            I => \Clock12MHz_c\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_8_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_8_4_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visibley_cry_7,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un21_beamy_cry_8,
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_4_0_\
        );

    \IN_MUX_bfv_12_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_5_0_\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_7_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_1_0_\
        );

    \IN_MUX_bfv_7_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_2_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2252\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2485\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_1_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNI0365_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2303\,
            in2 => \_gnd_net_\,
            in3 => \N__2291\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4_c_RNIZ0Z0365\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPF3_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2309\,
            in2 => \N__4052\,
            in3 => \N__2288\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5_c_RNIOPFZ0Z3\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6_c_RNIBRH7_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__2443\,
            in1 => \N__2264\,
            in2 => \N__2276\,
            in3 => \N__2285\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_axb_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2282\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23\,
            ltout => \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2SZ0Z23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un47_sum_cry_7_c_RNI2S23_0_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2279\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3U_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2262\,
            in2 => \_gnd_net_\,
            in3 => \N__2263\,
            lcout => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIG3UZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2467\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_2_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2267\,
            lcout => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1F_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2312\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un40_sum_cry_4_c_RNIO1FZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2468\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un40_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIS9H2_9_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__2847\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2917\,
            lcout => \N_132\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2T15_1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__3096\,
            in1 => \N__3133\,
            in2 => \N__3050\,
            in3 => \N__2730\,
            lcout => OPEN,
            ltout => \un5_beamx_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIP1J7_5_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2963\,
            in2 => \N__2297\,
            in3 => \N__3004\,
            lcout => OPEN,
            ltout => \un5_beamx_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI9DLC_0_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2885\,
            in1 => \N__2588\,
            in2 => \N__2294\,
            in3 => \N__2765\,
            lcout => un5_beamx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__2347\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4272\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4179\,
            ce => \N__3548\,
            sr => \_gnd_net_\
        );

    \beamY_0_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2346\,
            in2 => \_gnd_net_\,
            in3 => \N__2769\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4179\,
            ce => \N__3548\,
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2731\,
            in2 => \N__2771\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => un21_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_2_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3131\,
            in2 => \_gnd_net_\,
            in3 => \N__2375\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => un21_beamy_cry_2,
            clk => \N__4178\,
            ce => \N__3543\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2348\,
            in1 => \N__3088\,
            in2 => \_gnd_net_\,
            in3 => \N__2372\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \N__4178\,
            ce => \N__3543\,
            sr => \_gnd_net_\
        );

    \beamY_4_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2354\,
            in1 => \N__3044\,
            in2 => \_gnd_net_\,
            in3 => \N__2369\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \N__4178\,
            ce => \N__3543\,
            sr => \_gnd_net_\
        );

    \beamY_5_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3002\,
            in2 => \_gnd_net_\,
            in3 => \N__2366\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \N__4178\,
            ce => \N__3543\,
            sr => \_gnd_net_\
        );

    \beamY_6_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2953\,
            in2 => \_gnd_net_\,
            in3 => \N__2363\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \N__4178\,
            ce => \N__3543\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__2349\,
            in1 => \N__2915\,
            in2 => \_gnd_net_\,
            in3 => \N__2360\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \N__4178\,
            ce => \N__3543\,
            sr => \_gnd_net_\
        );

    \beamY_8_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2881\,
            in2 => \_gnd_net_\,
            in3 => \N__2357\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \N__4178\,
            ce => \N__3543\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__2846\,
            in1 => \N__2353\,
            in2 => \_gnd_net_\,
            in3 => \N__2315\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4177\,
            ce => \N__3544\,
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3170\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FE_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2419\,
            in2 => \N__2387\,
            in3 => \N__2447\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4_c_RNIU4FEZ0\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HH_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2444\,
            in2 => \N__2432\,
            in3 => \N__2423\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5_c_RNI00HHZ0\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6_c_RNI4PN01_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3226\,
            in1 => \N__2420\,
            in2 => \N__2411\,
            in3 => \N__2402\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2399\,
            in2 => \_gnd_net_\,
            in3 => \N__2393\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0\,
            ltout => \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SGZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un54_sum_cry_7_c_RNIB0SG_0_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2390\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2486\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3489\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3421\,
            in2 => \_gnd_net_\,
            in3 => \N__2378\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3454\,
            in2 => \N__4056\,
            in3 => \N__2492\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2690\,
            in2 => \_gnd_net_\,
            in3 => \N__2489\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2669\,
            in2 => \N__4057\,
            in3 => \N__2474\,
            lcout => \un1_beamX_if_generate_plus_mult1_un47_sum\,
            ltout => OPEN,
            carryin => un5_visiblex_cry_7,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2648\,
            in2 => \_gnd_net_\,
            in3 => \N__2471\,
            lcout => \un1_beamX_if_generate_plus_mult1_un40_sum\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2510\,
            in2 => \N__2531\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2545\,
            in2 => \_gnd_net_\,
            in3 => \N__2459\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__4182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3393\,
            in2 => \_gnd_net_\,
            in3 => \N__2456\,
            lcout => \N_97\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__4182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3536\,
            in1 => \N__3496\,
            in2 => \_gnd_net_\,
            in3 => \N__2453\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__4182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3427\,
            in2 => \_gnd_net_\,
            in3 => \N__2450\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__4182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3459\,
            in2 => \_gnd_net_\,
            in3 => \N__2561\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__4182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2693\,
            in2 => \_gnd_net_\,
            in3 => \N__2558\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__4182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2672\,
            in2 => \_gnd_net_\,
            in3 => \N__2555\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__4182\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2647\,
            in2 => \_gnd_net_\,
            in3 => \N__2552\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_4_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__4181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__3687\,
            in1 => \N__3523\,
            in2 => \_gnd_net_\,
            in3 => \N__2549\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNITFL_1_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2523\,
            in1 => \N__2507\,
            in2 => \N__2546\,
            in3 => \N__3458\,
            lcout => un3_beamx_i_i_a2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__2509\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2524\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__3524\,
            in1 => \N__2508\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4181\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNINLG_7_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__2644\,
            in1 => \N__2670\,
            in2 => \_gnd_net_\,
            in3 => \N__2691\,
            lcout => \N_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_15_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000011"
        )
    port map (
            in0 => \N__2692\,
            in1 => \N__2671\,
            in2 => \N__3461\,
            in3 => \N__2645\,
            lcout => OPEN,
            ltout => \Pixel_0_sqmuxa_i_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_14_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101001011000"
        )
    port map (
            in0 => \N__2646\,
            in1 => \N__3422\,
            in2 => \N__2624\,
            in3 => \N__3493\,
            lcout => \Pixel_0_sqmuxa_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQUP3_9_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__2849\,
            in1 => \N__2884\,
            in2 => \_gnd_net_\,
            in3 => \N__2918\,
            lcout => un1_beamylto9_0_a2_1,
            ltout => \un1_beamylto9_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSync_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__2782\,
            in1 => \N__3143\,
            in2 => \N__2621\,
            in3 => \N__2729\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_11_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__3141\,
            in1 => \N__2727\,
            in2 => \N__3097\,
            in3 => \N__2763\,
            lcout => OPEN,
            ltout => \N_84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_8_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010001"
        )
    port map (
            in0 => \N__2962\,
            in1 => \N__3005\,
            in2 => \N__2591\,
            in3 => \N__3049\,
            lcout => \N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_13_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__3705\,
            in1 => \N__2848\,
            in2 => \N__3689\,
            in3 => \N__2883\,
            lcout => \Pixel_0_sqmuxa_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_12_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__2764\,
            in1 => \N__3142\,
            in2 => \N__2783\,
            in3 => \N__2728\,
            lcout => OPEN,
            ltout => \N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_9_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__2587\,
            in1 => \N__2576\,
            in2 => \N__2570\,
            in3 => \N__2567\,
            lcout => OPEN,
            ltout => \Pixel_0_sqmuxa_i_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2810\,
            in2 => \N__2804\,
            in3 => \N__2801\,
            lcout => \Pixel_0_sqmuxa_i_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3969\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PP_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3882\,
            in1 => \N__3971\,
            in2 => \_gnd_net_\,
            in3 => \N__2795\,
            lcout => \un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0_c_RNIQ0PPZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un26_sum_cry_3_s0,
            carryout => un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0_c_RNIR53K_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3883\,
            in1 => \N__3970\,
            in2 => \_gnd_net_\,
            in3 => \N__2792\,
            lcout => un1_visibley_if_generate_plus_mult1_un33_sum_axb_6,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un26_sum_cry_4_s0,
            carryout => un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3884\,
            in2 => \N__3893\,
            in3 => \N__2789\,
            lcout => \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0\,
            ltout => \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCKZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un26_sum_cry_5_s0_c_RNIICCK_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2786\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un33_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIA525_3_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2995\,
            in1 => \N__3037\,
            in2 => \N__3098\,
            in3 => \N__2961\,
            lcout => \N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_0_c_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2770\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => un5_visibley_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_0_c_RNIJVSB_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2732\,
            in3 => \N__2696\,
            lcout => \un5_visibley_cry_0_c_RNIJVSBZ0\,
            ltout => OPEN,
            carryin => un5_visibley_cry_0,
            carryout => un5_visibley_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_1_c_RNIL2UB_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4000\,
            in2 => \N__3132\,
            in3 => \N__3101\,
            lcout => un1_visibley_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_1,
            carryout => un5_visibley_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_2_c_RNIN5VB_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3089\,
            in3 => \N__3053\,
            lcout => un1_visibley_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_2,
            carryout => un5_visibley_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_3_c_RNIP80C_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4001\,
            in2 => \N__3045\,
            in3 => \N__3008\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_3,
            carryout => un5_visibley_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_4_c_RNIRB1C_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3003\,
            in3 => \N__2966\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_4,
            carryout => un5_visibley_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_5_c_RNITE2C_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4002\,
            in2 => \N__2954\,
            in3 => \N__2921\,
            lcout => un1_visibley_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_5,
            carryout => un5_visibley_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_6_c_RNIVH3C_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4031\,
            in2 => \N__2916\,
            in3 => \N__2888\,
            lcout => un1_visibley_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => un5_visibley_cry_6,
            carryout => un5_visibley_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_7_c_RNI1L4C_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4035\,
            in2 => \N__2882\,
            in3 => \N__2852\,
            lcout => un1_visibley_if_generate_plus_mult1_un33_sum,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => un5_visibley_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_8_c_RNI3O5C_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2836\,
            in2 => \_gnd_net_\,
            in3 => \N__2813\,
            lcout => un1_visibley_if_generate_plus_mult1_un26_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3316\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FE21_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3202\,
            in2 => \N__3155\,
            in3 => \N__3230\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4_c_RNI3FEZ0Z21\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQE1_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3227\,
            in2 => \N__3215\,
            in3 => \N__3206\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5_c_RNI5FQEZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6_c_RNIAJ623_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3370\,
            in1 => \N__3203\,
            in2 => \N__3194\,
            in3 => \N__3185\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3182\,
            in2 => \_gnd_net_\,
            in3 => \N__3176\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1\,
            ltout => \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279GZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un61_sum_cry_7_c_RNI279G1_0_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3173\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3169\,
            lcout => \un1_beamX_if_generate_plus_mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3295\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BK1_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3346\,
            in2 => \N__3305\,
            in3 => \N__3146\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4_c_RNIV6BKZ0Z1\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNK2_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3371\,
            in2 => \N__3359\,
            in3 => \N__3350\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5_c_RNI8KNKZ0Z2\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6_c_RNIQBD56_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3256\,
            in1 => \N__3347\,
            in2 => \N__3338\,
            in3 => \N__3329\,
            lcout => \un1_beamX_if_generate_plus_mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFL843_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3326\,
            in2 => \_gnd_net_\,
            in3 => \N__3320\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_cry_7_c_RNIFLZ0Z843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3317\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3296\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3585\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58A_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3238\,
            in2 => \N__3287\,
            in3 => \N__3278\,
            lcout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_RNIP58AZ0\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_7_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3275\,
            in2 => \N__3257\,
            in3 => \N__3269\,
            lcout => \Pixel_1_RNOZ0Z_7\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_5\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3239\,
            in2 => \N__3266\,
            in3 => \N__3252\,
            lcout => \un1_beamX_if_generate_plus_mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_6\,
            carryout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMD6_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3605\,
            in2 => \_gnd_net_\,
            in3 => \N__3599\,
            lcout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6\,
            ltout => \un1_beamX_if_generate_plus_mult1_un75_sum_cry_7_c_RNITMMDZ0Z6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_2_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111110110000"
        )
    port map (
            in0 => \N__3586\,
            in1 => \N__3575\,
            in2 => \N__3596\,
            in3 => \N__3593\,
            lcout => \N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_beamX_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__4053\,
            in1 => \N__3587\,
            in2 => \_gnd_net_\,
            in3 => \N__3497\,
            lcout => un5_visiblex_i,
            ltout => \un5_visiblex_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_1_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110101110011"
        )
    port map (
            in0 => \N__3398\,
            in1 => \N__3574\,
            in2 => \N__3566\,
            in3 => \N__3563\,
            lcout => \N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_10_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4150\,
            in2 => \_gnd_net_\,
            in3 => \N__4273\,
            lcout => \G_7_0_a4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNIHUU5_10_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__3686\,
            in1 => \N__3423\,
            in2 => \N__3397\,
            in3 => \N__3494\,
            lcout => OPEN,
            ltout => \un3_beamx_i_i_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_RNI5457_1_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3557\,
            in2 => \N__3551\,
            in3 => \N__3706\,
            lcout => \beamX_RNI5457Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_RNO_0_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3495\,
            in1 => \N__3460\,
            in2 => \N__3428\,
            in3 => \N__3392\,
            lcout => OPEN,
            ltout => \N_130_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSync_1_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__3707\,
            in1 => \_gnd_net_\,
            in2 => \N__3692\,
            in3 => \N__3688\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3616\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJI2_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3753\,
            in2 => \N__3716\,
            in3 => \N__3635\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_RNIIPJIZ0Z2\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6P3_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3833\,
            in2 => \N__3758\,
            in3 => \N__3632\,
            lcout => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_3_c_RNINV6PZ0Z3\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QOR3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3757\,
            in2 => \N__3824\,
            in3 => \N__3629\,
            lcout => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_4_c_RNI7QORZ0Z3\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_5_c_RNIEFE58_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4339\,
            in1 => \N__3812\,
            in2 => \N__3734\,
            in3 => \N__3626\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3794\,
            in2 => \_gnd_net_\,
            in3 => \N__3623\,
            lcout => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94\,
            ltout => \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FIZ0Z94_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_cry_6_c_RNI4FI94_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3620\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un47_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un47_sum_sbtinv_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3617\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3724\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVF1_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3839\,
            in2 => \N__3783\,
            in3 => \N__3827\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_2_c_RNI9AVFZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GI1_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3776\,
            in2 => \N__4088\,
            in3 => \N__3815\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_3_c_RNIO2GIZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6II1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4076\,
            in2 => \N__3784\,
            in3 => \N__3806\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_4_c_RNIQ6IIZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_5_c_RNI9GRQ3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3752\,
            in1 => \N__3935\,
            in2 => \N__3803\,
            in3 => \N__3788\,
            lcout => un1_visibley_if_generate_plus_mult1_un47_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__3922\,
            in1 => \N__3908\,
            in2 => \N__3785\,
            in3 => \N__3761\,
            lcout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1\,
            ltout => \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMSJQ1_0_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3737\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3847\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0I_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4036\,
            in2 => \N__3857\,
            in3 => \N__4079\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_2_c_RNILH0IZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1I_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3873\,
            in2 => \N__4054\,
            in3 => \N__4070\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_3_c_RNIMJ1IZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULV_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4067\,
            in2 => \N__4055\,
            in3 => \N__3926\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_4_c_RNIEULVZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un33_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3923\,
            in3 => \N__3899\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un33_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un33_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_LUT4_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3896\,
            lcout => \un1_visibley_if_generate_plus_mult1_un33_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visibley_cry_8_c_RNI3O5C_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3872\,
            lcout => \un5_visibley_cry_8_c_RNI3O5CZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un33_sum_sbtinv_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3848\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un33_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_4_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__4417\,
            in1 => \N__4402\,
            in2 => \N__4154\,
            in3 => \N__4094\,
            lcout => OPEN,
            ltout => \N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_0_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001011"
        )
    port map (
            in0 => \N__4277\,
            in1 => \N__4115\,
            in2 => \N__4253\,
            in3 => \N__4391\,
            lcout => OPEN,
            ltout => \N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000000101"
        )
    port map (
            in0 => \N__4250\,
            in1 => \N__4238\,
            in2 => \N__4229\,
            in3 => \N__4226\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4149\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTP21_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4385\,
            in2 => \N__4462\,
            in3 => \N__4121\,
            lcout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_2_c_RNILGTPZ0Z21\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78K1_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4457\,
            in2 => \N__4508\,
            in3 => \N__4118\,
            lcout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_3_c_RNIAP78KZ0Z1\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_6_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4496\,
            in2 => \N__4463\,
            in3 => \N__4109\,
            lcout => \Pixel_1_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4487\,
            in2 => \N__4106\,
            in3 => \N__4453\,
            lcout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_invZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMI32_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4478\,
            in3 => \N__4097\,
            lcout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32\,
            ltout => \un1_visibley_if_generate_plus_mult1_un75_sum_cry_6_c_RNIGAMIZ0Z32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_1_RNO_5_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4427\,
            in1 => \N__4418\,
            in2 => \N__4406\,
            in3 => \N__4403\,
            lcout => \N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_sbtinv_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4526\,
            lcout => un1_visibley_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4540\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TM4_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4347\,
            in2 => \N__4379\,
            in3 => \N__4367\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_2_c_RNI52TMZ0Z4\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICA117_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4364\,
            in2 => \N__4352\,
            in3 => \N__4355\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_3_c_RNICAZ0Z117\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIIL78_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4351\,
            in2 => \N__4328\,
            in3 => \N__4316\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIILZ0Z78\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_5_c_RNIA6LKG_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4643\,
            in1 => \N__4313\,
            in2 => \N__4304\,
            in3 => \N__4292\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4289\,
            in2 => \_gnd_net_\,
            in3 => \N__4280\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8\,
            ltout => \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCAZ0Z8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_cry_6_c_RNI7NCA8_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4544\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4541\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4525\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPH_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4572\,
            in2 => \N__4436\,
            in3 => \N__4499\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_RNI3TLPHZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85Q_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4676\,
            in2 => \N__4577\,
            in3 => \N__4490\,
            lcout => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_3_c_RNI0K85QZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPU_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4576\,
            in2 => \N__4661\,
            in3 => \N__4481\,
            lcout => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_4_c_RNITRQPUZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_5_c_RNIKSOE32_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4461\,
            in1 => \N__4619\,
            in2 => \N__4553\,
            in3 => \N__4469\,
            lcout => un1_visibley_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNA21_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4595\,
            in2 => \_gnd_net_\,
            in3 => \N__4466\,
            lcout => \un1_visibley_if_generate_plus_mult1_un68_sum_cry_6_c_RNIEKNAZ0Z21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_sbtinv_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4709\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4708\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_5_0_\,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQN8_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4644\,
            in2 => \N__4685\,
            in3 => \N__4670\,
            lcout => \un1_visibley_if_generate_plus_mult1_un54_sum_sbtinv_RNI4UQNZ0Z8\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCD_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4667\,
            in2 => \N__4649\,
            in3 => \N__4652\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_3_c_RNI04CCDZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMF_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4648\,
            in2 => \N__4628\,
            in3 => \N__4613\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_4_c_RNI8EHMFZ0\,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_5_c_RNIGF1T11_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__4571\,
            in1 => \N__4610\,
            in2 => \N__4604\,
            in3 => \N__4589\,
            lcout => un1_visibley_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => un1_visibley_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => un1_visibley_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4586\,
            in2 => \_gnd_net_\,
            in3 => \N__4580\,
            lcout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0\,
            ltout => \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVGZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un1_visibley_if_generate_plus_mult1_un61_sum_cry_6_c_RNI1NQVG_0_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4556\,
            in3 => \_gnd_net_\,
            lcout => un1_visibley_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
