-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2014.12.27052

-- Build Date:         Dec  8 2014 15:16:02

-- File Generated:     Jun 24 2015 00:16:13

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "SimpleVGA" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of SimpleVGA
entity SimpleVGA is
port (
    VSync : out std_logic;
    SDATA : in std_logic;
    SCLK1 : out std_logic;
    Pixel : out std_logic;
    HSync : out std_logic;
    nCS2 : out std_logic;
    SCLK2 : out std_logic;
    Clock12MHz : in std_logic;
    nCS1 : out std_logic);
end SimpleVGA;

-- Architecture of SimpleVGA
-- View name is \INTERFACE\
architecture \INTERFACE\ of SimpleVGA is

signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16024\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15499\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15205\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15085\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15065\ : std_logic;
signal \N__15062\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14782\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14491\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14455\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13715\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13607\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \Clock50MHz.PixelClock\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal un21_beamy_cry_1 : std_logic;
signal un21_beamy_cry_2 : std_logic;
signal un21_beamy_cry_3 : std_logic;
signal un21_beamy_cry_4 : std_logic;
signal un21_beamy_cry_5 : std_logic;
signal un21_beamy_cry_6 : std_logic;
signal un21_beamy_cry_7 : std_logic;
signal un21_beamy_cry_8 : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOGZ0Z53\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOSZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRSZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LKZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01_cascade_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0 : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOLZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IGZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMGZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0 : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICMZ0Z321\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPMZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KHZ0Z2\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0 : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CRZ0Z2\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGIZ0Z3\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJZ0Z6874\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7 : std_logic;
signal \un21_beamy_cry_4_c_RNIGUAZ0Z3\ : std_logic;
signal \un21_beamy_cry_6_c_RNIK4DZ0Z3\ : std_logic;
signal \beamY_fastZ0Z_7\ : std_logic;
signal \beamY_fastZ0Z_5\ : std_logic;
signal \un21_beamy_cry_1_c_RNIALZ0Z73\ : std_logic;
signal un5_visibley_c6_0_0_0 : std_logic;
signal \beamY_fast_RNI35GAZ0Z_2_cascade_\ : std_logic;
signal \un21_beamy_cry_2_c_RNICOZ0Z83\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2LZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RCZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5 : std_logic;
signal \beamY_RNIFJ0L_0Z0Z_8\ : std_logic;
signal \beamY_RNI19IJ_0Z0Z_9\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7 : std_logic;
signal \beamY_i_2_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__chessboardpixel_un200_pixellto4Z0Z_1_cascade_\ : std_logic;
signal \chessboardpixel_un200_pixellt10_cascade_\ : std_logic;
signal \chessboardpixel_un200_pixel_0_1_cascade_\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5 : std_logic;
signal \beamY_i_2\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81BZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEGZ0Z5\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODGZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87VZ0Z68\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4JZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05UZ0Z8\ : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGKZ0\ : std_logic;
signal chessboardpixel_un174_pixel_0_1 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0 : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHFZ0\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJZ0Z5\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0\ : std_logic;
signal \un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1Z0Z_1\ : std_logic;
signal \un114_pixel_1_0_3__un1_beamylto9Z0Z_0_cascade_\ : std_logic;
signal \un4_beamylt6_cascade_\ : std_logic;
signal un5_visibley_ac0_11_d : std_logic;
signal un5_visibley_ac0_11_0_1 : std_logic;
signal \un114_pixel_1_0_3__un1_beamylto9_3\ : std_logic;
signal \beamY_fastZ0Z_2\ : std_logic;
signal \beamYZ0Z_5\ : std_logic;
signal \beamY_fastZ0Z_3\ : std_logic;
signal \beamY_fast_RNIM4P7Z0Z_2_cascade_\ : std_logic;
signal \beamYZ0Z_6\ : std_logic;
signal un5_visibley_c5 : std_logic;
signal \un5_visibley_c5_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__un5_beamxZ0Z_5_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__g0_1Z0Z_0_cascade_\ : std_logic;
signal un4_beamylt8_0 : std_logic;
signal un5_visibley_c2 : std_logic;
signal un1_beamy_4 : std_logic;
signal \beamYZ0Z_8\ : std_logic;
signal \beamYZ0Z_9\ : std_logic;
signal \un114_pixel_1_0_3__un8_beamylto9Z0Z_1_cascade_\ : std_logic;
signal \beamYZ0Z_7\ : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_cZ0Z4\ : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_cZ0Z4_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\ : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_\ : std_logic;
signal if_generate_plus_mult1_un68_sum_axbxc3 : std_logic;
signal \row_1_if_generate_plus_mult1_un68_sum_c5_0_nsZ0Z_1\ : std_logic;
signal row_1_if_generate_plus_mult1_un68_sum_c5 : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axbxc3 : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5_cascade_\ : std_logic;
signal row_1_if_generate_plus_mult1_un61_sum_c5 : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_c5_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0\ : std_logic;
signal if_generate_plus_mult1_un68_sum_c5_0_bm : std_logic;
signal row_1_if_generate_plus_mult1_un61_sum_ac0_7_c : std_logic;
signal \bfn_4_11_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KCZ0Z4\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGSZ0Z6\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8 : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal counter_cry_1 : std_logic;
signal counter_cry_2 : std_logic;
signal counter_cry_3 : std_logic;
signal counter_cry_4 : std_logic;
signal \slaveselect_1_0_4_cascade_\ : std_logic;
signal counter_30 : std_logic;
signal \un3_slaveselect_cascade_\ : std_logic;
signal counter_29 : std_logic;
signal \counter_31_cascade_\ : std_logic;
signal \counterZ0Z_0\ : std_logic;
signal \counterZ0Z_3\ : std_logic;
signal \counterZ0Z_1\ : std_logic;
signal \un1_counterlto3_0_cascade_\ : std_logic;
signal \counterZ0Z_2\ : std_logic;
signal \g0_0_1_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_c5 : std_logic;
signal un5_visibley_0_29 : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_c5_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_0_1_5 : std_logic;
signal \chary_if_generate_plus_mult1_un68_sum_c4_0_cascade_\ : std_logic;
signal g0_0_3 : std_logic;
signal \g1_0_cascade_\ : std_logic;
signal un4_beamylt6 : std_logic;
signal \chary_if_generate_plus_mult1_un75_sum_c5_N_9_cascade_\ : std_logic;
signal g0_1_2 : std_logic;
signal g0_2_0 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_1_0_1_0_3 : std_logic;
signal \beamY_RNINITP61Z0Z_5_cascade_\ : std_logic;
signal \beamY_RNINITP61_1Z0Z_5\ : std_logic;
signal chary_if_generate_plus_mult1_un40_sum_axb3 : std_logic;
signal \chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_axbxc5_2 : std_logic;
signal \chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un40_sum_c4 : std_logic;
signal chary_if_generate_plus_mult1_un47_sum_c5 : std_logic;
signal \beamY_RNITURI3_0Z0Z_7_cascade_\ : std_logic;
signal \beamY_RNITURI3Z0Z_7\ : std_logic;
signal un4_beamy_0 : std_logic;
signal un8_beamy : std_logic;
signal \un114_pixel_1_0_3__un15_beamyZ0Z_2\ : std_logic;
signal \un1_beamx_2_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__un5_beamxZ0Z_3\ : std_logic;
signal \beamYZ0Z_4\ : std_logic;
signal \un114_pixel_1_0_3__g0_1Z0Z_3\ : std_logic;
signal \un114_pixel_1_0_3__un18_beamylto9Z0Z_2_cascade_\ : std_logic;
signal un18_beamylt10_0 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum : std_logic;
signal un13_beamylt7 : std_logic;
signal if_generate_plus_mult1_un75_sum_axbxc5 : std_logic;
signal if_generate_plus_mult1_un75_sum_axbxc3 : std_logic;
signal \row_1_if_generate_plus_mult1_un82_sum_axb4_i_cascade_\ : std_logic;
signal \row_1_if_generate_plus_mult1_un82_sum_ac0_7_0Z0Z_1\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal un8_beamx_cry_1 : std_logic;
signal un8_beamx_cry_2 : std_logic;
signal un8_beamx_cry_3 : std_logic;
signal un8_beamx_cry_4 : std_logic;
signal un8_beamx_cry_5 : std_logic;
signal un8_beamx_cry_6 : std_logic;
signal un8_beamx_cry_7 : std_logic;
signal un8_beamx_cry_8 : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal un8_beamx_cry_9 : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un19_sum_cry_2 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i : std_logic;
signal counter_27 : std_logic;
signal \counterZ0Z_5\ : std_logic;
signal slaveselect_1_0_4 : std_logic;
signal un1_slaveselect_1_i : std_logic;
signal un3_slaveselect : std_logic;
signal counter_28 : std_logic;
signal \counterZ0Z_4\ : std_logic;
signal \slaveselectZ0\ : std_logic;
signal un1_counter_0 : std_logic;
signal \nCS1_c\ : std_logic;
signal \nCS1_0_sqmuxa\ : std_logic;
signal \beamY_RNI2TEJF4Z0Z_4_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__g0_8Z0Z_1\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_0_3_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__g0_1Z0Z_1_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_0_3 : std_logic;
signal \un114_pixel_1_0_3__g0_3Z0Z_0_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un75_sum_i_0_5 : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c4_0 : std_logic;
signal \un114_pixel_1_0_3__g0Z0Z_1_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_0_0_0_0_5 : std_logic;
signal g2 : std_logic;
signal \un114_pixel_1_0_3__g0Z0Z_3_cascade_\ : std_logic;
signal \beamY_RNITFRN03Z0Z_5\ : std_logic;
signal chary_if_generate_plus_mult1_un75_sum_c5 : std_logic;
signal \beamY_RNIH9THADZ0Z_4_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb3_0 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_7_d : std_logic;
signal \beamY_RNIKHPCA1Z0Z_4\ : std_logic;
signal \chary_if_generate_plus_mult1_un61_sum_ac0_7_d_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_axb4 : std_logic;
signal \beamY_RNI2TEJF4Z0Z_4\ : std_logic;
signal chary_if_generate_plus_mult1_un68_sum_c4 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb4_0 : std_logic;
signal \g0_0_x2_1_1_cascade_\ : std_logic;
signal g0_3_2 : std_logic;
signal \beamY_RNIARUFBZ0Z_5_cascade_\ : std_logic;
signal \beamY_RNIGS0LBZ0Z_5\ : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_c5 : std_logic;
signal \chary_if_generate_plus_mult1_un54_sum_c5_cascade_\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0 : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axb3_0_0 : std_logic;
signal \beamY_RNIDO3IZ0Z_9\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0 : std_logic;
signal g0_4_2 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_axb3 : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum : std_logic;
signal chary_if_generate_plus_mult1_un54_sum_axbxc5_1 : std_logic;
signal \beamY_RNI2MTA1Z0Z_9\ : std_logic;
signal \chary_if_generate_plus_mult1_un54_sum_c4_cascade_\ : std_logic;
signal \beamY_RNICG8P9Z0Z_7\ : std_logic;
signal chary_if_generate_plus_mult1_un61_sum_axbxc5_1 : std_logic;
signal \un3_beamx_0_cascade_\ : std_logic;
signal un1_beamx_2 : std_logic;
signal \HSync_c\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_1 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8VZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_cry_4 : std_logic;
signal un1_beamxlt10_0 : std_logic;
signal \beamXZ0Z_10\ : std_logic;
signal \un114_pixel_1_0_3__un3_beamxZ0Z_5_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__un3_beamxZ0Z_7\ : std_logic;
signal un18_beamylt4 : std_logic;
signal \charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO\ : std_logic;
signal \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKFZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un19_sum_i : std_logic;
signal \bfn_6_10_0_\ : std_logic;
signal \beamXZ0Z_1\ : std_logic;
signal un5_visiblex_cry_0 : std_logic;
signal \beamXZ0Z_2\ : std_logic;
signal un5_visiblex_cry_1 : std_logic;
signal \beamXZ0Z_3\ : std_logic;
signal un5_visiblex_cry_2 : std_logic;
signal \beamXZ0Z_4\ : std_logic;
signal un5_visiblex_cry_3 : std_logic;
signal \beamXZ0Z_5\ : std_logic;
signal un5_visiblex_cry_4 : std_logic;
signal \beamXZ0Z_6\ : std_logic;
signal un5_visiblex_cry_5 : std_logic;
signal \beamXZ0Z_7\ : std_logic;
signal un5_visiblex_cry_6 : std_logic;
signal un5_visiblex_cry_7 : std_logic;
signal \beamXZ0Z_8\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \beamXZ0Z_9\ : std_logic;
signal un5_visiblex_cry_8 : std_logic;
signal \un116_pixel_3_bm_2_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__N_5_1_0\ : std_logic;
signal \un114_pixel_1_0_3__un116_pixel_4_ns_1_0_7_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__g2_1Z0Z_0\ : std_logic;
signal \beamY_RNIH9THADZ0Z_4\ : std_logic;
signal \beamYZ0Z_3\ : std_logic;
signal \N_345_0_0_1\ : std_logic;
signal \font_un28_pixel_29_cascade_\ : std_logic;
signal \un116_pixel_5_am_6_cascade_\ : std_logic;
signal g1_1 : std_logic;
signal g0_0_x2_1 : std_logic;
signal \un114_pixel_1_0_3__un116_pixel_2_ns_1Z0Z_2_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__un116_pixel_5_ns_1Z0Z_2_cascade_\ : std_logic;
signal \un116_pixel_5_ns_1Z0Z_4_cascade_\ : std_logic;
signal un116_pixel_5_ns_2 : std_logic;
signal \N_362\ : std_logic;
signal \un116_pixel_7_ns_1_6_cascade_\ : std_logic;
signal \N_379\ : std_logic;
signal un116_pixel_3_ns_2 : std_logic;
signal \beamY_RNI57H3N31_0Z0Z_1_cascade_\ : std_logic;
signal \beamY_RNI896FQ3Z0Z_0\ : std_logic;
signal \beamY_RNI896FQ3Z0Z_0_cascade_\ : std_logic;
signal \beamY_RNI57H3N31Z0Z_1\ : std_logic;
signal \un116_pixel_2_ns_1_0_6_cascade_\ : std_logic;
signal \beamY_RNIGO5PPVZ0Z_0\ : std_logic;
signal \N_41\ : std_logic;
signal un3_beamx_0 : std_logic;
signal un5_beamx_0 : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_iZ0\ : std_logic;
signal \row_1_if_generate_plus_mult1_un54_sum_cZ0Z5\ : std_logic;
signal un5_rowlto3_i : std_logic;
signal \bfn_7_8_0_\ : std_logic;
signal \N_575_i\ : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un61_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal \bfn_7_9_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HLZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\ : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_i_5 : std_logic;
signal \bfn_7_10_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072\ : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_cry_4 : std_logic;
signal charx_if_generate_plus_mult1_un33_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un26_sum_i : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_2 : std_logic;
signal \N_204_0_i\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_0_cry_4 : std_logic;
signal un5_visiblex_i_25 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_cry_3_ma : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un54_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_4_l_fx : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3\ : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEBZ0Z2\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLITZ0Z2\ : std_logic;
signal charx_if_generate_plus_mult1_un40_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6\ : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0OZ0Z3\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCDZ0Z16\ : std_logic;
signal charx_if_generate_plus_mult1_un47_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal charx_if_generate_plus_mult1_un54_sum : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLMZ0Z67\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSAZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0_cascade_\ : std_logic;
signal \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un54_sum_i_5 : std_logic;
signal \VSync_c\ : std_logic;
signal un116_pixel_3_am_2 : std_logic;
signal \N_1556_0_cascade_\ : std_logic;
signal \N_347_0\ : std_logic;
signal font_un28_pixel_0_29 : std_logic;
signal \N_368_0\ : std_logic;
signal \un114_pixel_1_0_3__font_un126_pixel_1_d_ns_1_0_cascade_\ : std_logic;
signal \N_389_0\ : std_logic;
signal \N_346_0_0_1\ : std_logic;
signal \g0_cascade_\ : std_logic;
signal \N_36_cascade_\ : std_logic;
signal \un116_pixel_3_ns_1_1_cascade_\ : std_logic;
signal \font_un3_pixel_29_cascade_\ : std_logic;
signal un116_pixel_5_bm_6 : std_logic;
signal un116_pixel_4_bm_1 : std_logic;
signal \beamY_RNI1C50FS3Z0Z_0_cascade_\ : std_logic;
signal \un116_pixel_3_bm_1_6_cascade_\ : std_logic;
signal \beamY_RNIOHI2NGZ0Z_0\ : std_logic;
signal \N_364_cascade_\ : std_logic;
signal \un116_pixel_7_ns_1_4_cascade_\ : std_logic;
signal \beamY_RNI2L0T663Z0Z_0\ : std_logic;
signal column_0111_1_0 : std_logic;
signal \beamY_RNI1J75181Z0Z_1\ : std_logic;
signal \font_un126_pixel_6_am_cascade_\ : std_logic;
signal un1_beamy_0 : std_logic;
signal \N_1075_0_cascade_\ : std_logic;
signal \N_400\ : std_logic;
signal \Pixel_r_rn_0_cascade_\ : std_logic;
signal \Pixel_c\ : std_logic;
signal \PixelClock_g\ : std_logic;
signal font_un28_pixel_0_0_29 : std_logic;
signal font_un126_pixel_2_bm : std_logic;
signal \un114_pixel_1_0_3__font_un126_pixel_7_d_ns_1_0_0\ : std_logic;
signal \beamY_RNIHHB5F01Z0Z_4\ : std_logic;
signal \beamYZ0Z_2\ : std_logic;
signal \beamY_RNI7OE17CZ0Z_0\ : std_logic;
signal \beamY_RNIVU1O9RZ0Z_1\ : std_logic;
signal font_un126_pixel_6_bm : std_logic;
signal \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\ : std_logic;
signal un15_beamy : std_logic;
signal \r_i1_mux_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_1_cascade_\ : std_logic;
signal chary_24 : std_logic;
signal \un114_pixel_1_0_3__font_un126_pixel_m_1_0_cascade_\ : std_logic;
signal chary_23 : std_logic;
signal \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3\ : std_logic;
signal un1_beamylto9 : std_logic;
signal \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3_cascade_\ : std_logic;
signal \Pixel_r_sn\ : std_logic;
signal \beamXZ0Z_0\ : std_logic;
signal \un114_pixel_1_0_3__font_un57_pixelZ0Z_0\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum : std_logic;
signal if_generate_plus_mult1_un61_sum_axbxc5 : std_logic;
signal \un114_pixel_1_0_3__un4_row_8Z0Z_3_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__un4_row_8_7Z0Z_1\ : std_logic;
signal chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum : std_logic;
signal chary_if_generate_plus_mult1_un33_sum_axb3 : std_logic;
signal if_generate_plus_mult1_un54_sum_s_5 : std_logic;
signal \un114_pixel_1_0_3__un4_row_8Z0Z_2\ : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_cZ0Z5\ : std_logic;
signal if_generate_plus_mult1_un68_sum_axbxc5 : std_logic;
signal \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2\ : std_logic;
signal \un114_pixel_1_0_3__un4_row_8Z0Z_7\ : std_logic;
signal \un114_pixel_1_0_3__un4_rowZ0Z_8\ : std_logic;
signal \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1\ : std_logic;
signal row_1_if_generate_plus_mult1_un82_sum_c5 : std_logic;
signal \un114_pixel_1_0_3__un4_rowZ0Z_8_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__Pixel_3_sqmuxaZ0Z_0\ : std_logic;
signal \Pixel_3_sqmuxa\ : std_logic;
signal \bfn_8_10_0_\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_4_c_invZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843_cascade_\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i : std_logic;
signal \un114_pixel_1_0_3__un4_row_8Z0Z_0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_i_5 : std_logic;
signal if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axb_2_sxZ0_cascade_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2_cascade_\ : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_2_l_fx : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_4 : std_logic;
signal \if_generate_plus_mult1_un47_sum_m_5_cascade_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_2 : std_logic;
signal if_generate_plus_mult1_un47_sum_m_5 : std_logic;
signal if_generate_plus_mult1_un54_sum_axb_3_l_fx : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum0_5 : std_logic;
signal \N_584_i\ : std_logic;
signal \N_37_i\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5RZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_1 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRDZ0\ : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BVZ0Z81\ : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_2 : std_logic;
signal \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0LZ0\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i_5 : std_logic;
signal charx_if_generate_plus_mult1_un75_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_3 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_axb_5 : std_logic;
signal charx_if_generate_plus_mult1_un68_sum_cry_4 : std_logic;
signal \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1\ : std_logic;
signal charx_if_generate_plus_mult1_un61_sum_i : std_logic;
signal \N_41_0\ : std_logic;
signal column_0111_0 : std_logic;
signal un116_pixel_3_ns_1_0_3 : std_logic;
signal \un114_pixel_1_0_3__g1Z0Z_4\ : std_logic;
signal \N_1583_0_cascade_\ : std_logic;
signal \N_26_0_0\ : std_logic;
signal \un116_pixel_2_amZ0Z_1_cascade_\ : std_logic;
signal un116_pixel_6_1 : std_logic;
signal \column_0001_0_cascade_\ : std_logic;
signal \beamY_RNILBST4T2Z0Z_1\ : std_logic;
signal \beamY_RNIT81CMJ2Z0Z_1_cascade_\ : std_logic;
signal font_un126_pixel_2_am : std_logic;
signal un116_pixel_4_am_1 : std_logic;
signal \N_36\ : std_logic;
signal \un116_pixel_5_amZ0Z_5\ : std_logic;
signal \un116_pixel_2_amZ0Z_5\ : std_logic;
signal \N_385\ : std_logic;
signal \N_325\ : std_logic;
signal \un116_pixel_2_bmZ0Z_1\ : std_logic;
signal \un114_pixel_1_0_3__un116_pixel_6_1Z0Z_1\ : std_logic;
signal un116_pixel_1_4 : std_logic;
signal \N_374_0\ : std_logic;
signal font_un3_pixel_29 : std_logic;
signal \un116_pixel_7_x0_0_cascade_\ : std_logic;
signal un116_pixel_7_x1_0 : std_logic;
signal un116_pixel_7_ns_0 : std_logic;
signal un116_pixel_2_bm_0 : std_logic;
signal \un114_pixel_1_0_3__un116_pixel_5_ns_1_0Z0Z_0\ : std_logic;
signal chessboardpixel_un152_pixel_24 : std_logic;
signal \un114_pixel_1_0_3__un116_pixel_6_1_1Z0Z_1\ : std_logic;
signal charx_if_generate_plus_mult1_un1_sum_axb1 : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3EZ0Z987\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\ : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8TZ0Z77\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\ : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3 : std_logic;
signal font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4 : std_logic;
signal \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\ : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77Z0Z_0\ : std_logic;
signal charx_i_23 : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1\ : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2\ : std_logic;
signal \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843\ : std_logic;
signal charx_i_24 : std_logic;
signal \bfn_9_11_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUHZ0Z2\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIVZ0Z6153\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i : std_logic;
signal charx_if_generate_plus_mult1_un40_sum : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal un5_visiblex_i_0_25 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_2 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_1 : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx : std_logic;
signal \N_858_i\ : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_2 : std_logic;
signal if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_4 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum_1_cry_4 : std_logic;
signal column_1_if_generate_plus_mult1_un47_sum1_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8 : std_logic;
signal charx_if_generate_plus_mult1_un33_sum : std_logic;
signal \N_66\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5LZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7JZ0Z31\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i : std_logic;
signal \Clock12MHz_c_g\ : std_logic;
signal \GB_BUFFER_Clock12MHz_c_g_THRU_CO\ : std_logic;
signal \N_1557_0\ : std_logic;
signal \N_41_0_0_0\ : std_logic;
signal \N_563\ : std_logic;
signal \un116_pixel_5_bmZ0Z_5_cascade_\ : std_logic;
signal un116_pixel_6_ns_1_5 : std_logic;
signal \un116_pixel_2_bmZ0Z_5\ : std_logic;
signal \un114_pixel_7_1_7__N_9_cascade_\ : std_logic;
signal \un114_pixel_1_0_3__un116_pixel_3_ns_1Z0Z_0_cascade_\ : std_logic;
signal \un114_pixel_6_1_5__N_8\ : std_logic;
signal \N_371\ : std_logic;
signal \beamY_RNIJUCG3J3Z0Z_1\ : std_logic;
signal charx_if_generate_plus_mult1_un75_sum : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \G_345\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_1 : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_2 : std_logic;
signal \G_346\ : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_3 : std_logic;
signal column_1_if_generate_plus_mult1_un82_sum_cry_4 : std_logic;
signal \un5_rowlto0_cascade_\ : std_logic;
signal \un116_pixel_1_bmZ0Z_1\ : std_logic;
signal \beamYZ0Z_1\ : std_logic;
signal \un116_pixel_1_bmZ0Z_1_cascade_\ : std_logic;
signal \beamY_RNIV622TRZ0Z_1\ : std_logic;
signal un116_pixel_2_ns_1_4 : std_logic;
signal \beamYZ0Z_0\ : std_logic;
signal \beamY_RNIITCG3J3Z0Z_0\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \column_1_if_generate_plus_mult1_un68_sum_iZ0\ : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_2_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_1 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_2_s : std_logic;
signal if_generate_plus_mult1_un75_sum_cry_3_s : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_2 : std_logic;
signal \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_3 : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\ : std_logic;
signal column_1_if_generate_plus_mult1_un75_sum_cry_4 : std_logic;
signal un5_rowlto1 : std_logic;
signal un5_rowlto0 : std_logic;
signal \un5_rowlto1_cascade_\ : std_logic;
signal un5_rowlto3 : std_logic;
signal un116_pixel_2_am_0 : std_logic;
signal if_generate_plus_mult1_un68_sum_cry_3_s : std_logic;
signal if_generate_plus_mult1_un75_sum_axb_4_l_fx : std_logic;
signal un5_rowlto2 : std_logic;
signal un5_rowlto2_i : std_logic;
signal charx_if_generate_plus_mult1_un68_sum : std_logic;
signal \column_1_if_generate_plus_mult1_un75_sum_iZ0\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5 : std_logic;
signal charx_if_generate_plus_mult1_un26_sum : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHGZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6QZ0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6 : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7 : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\ : std_logic;
signal \CO3_0\ : std_logic;
signal chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\ : std_logic;
signal \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKNZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \Clock12MHz_wire\ : std_logic;
signal \VSync_wire\ : std_logic;
signal \HSync_wire\ : std_logic;
signal \nCS1_wire\ : std_logic;
signal \Pixel_wire\ : std_logic;
signal \nCS2_wire\ : std_logic;
signal \SCLK1_wire\ : std_logic;
signal \SCLK2_wire\ : std_logic;
signal \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \Clock12MHz_wire\ <= Clock12MHz;
    VSync <= \VSync_wire\;
    HSync <= \HSync_wire\;
    nCS1 <= \nCS1_wire\;
    Pixel <= \Pixel_wire\;
    nCS2 <= \nCS2_wire\;
    SCLK1 <= \SCLK1_wire\;
    SCLK2 <= \SCLK2_wire\;
    \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \Clock50MHz.PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \Clock50MHz.PixelClock\,
            REFERENCECLK => \N__14306\,
            RESETB => \N__16348\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \Clock50MHz.PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \Clock12MHz_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__16511\,
            GLOBALBUFFEROUTPUT => \Clock12MHz_c_g\
        );

    \Clock12MHz_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16513\,
            DIN => \N__16512\,
            DOUT => \N__16511\,
            PACKAGEPIN => \Clock12MHz_wire\
        );

    \Clock12MHz_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__16513\,
            PADOUT => \N__16512\,
            PADIN => \N__16511\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16502\,
            DIN => \N__16501\,
            DOUT => \N__16500\,
            PACKAGEPIN => \VSync_wire\
        );

    \VSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16502\,
            PADOUT => \N__16501\,
            PADIN => \N__16500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11668\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \HSync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16493\,
            DIN => \N__16492\,
            DOUT => \N__16491\,
            PACKAGEPIN => \HSync_wire\
        );

    \HSync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16493\,
            PADOUT => \N__16492\,
            PADIN => \N__16491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16484\,
            DIN => \N__16483\,
            DOUT => \N__16482\,
            PACKAGEPIN => \nCS1_wire\
        );

    \nCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16484\,
            PADOUT => \N__16483\,
            PADIN => \N__16482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8818\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Pixel_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16475\,
            DIN => \N__16474\,
            DOUT => \N__16473\,
            PACKAGEPIN => \Pixel_wire\
        );

    \Pixel_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16475\,
            PADOUT => \N__16474\,
            PADIN => \N__16473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11896\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCS2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16466\,
            DIN => \N__16465\,
            DOUT => \N__16464\,
            PACKAGEPIN => \nCS2_wire\
        );

    \nCS2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__16466\,
            PADOUT => \N__16465\,
            PADIN => \N__16464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8817\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCLK1_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16457\,
            DIN => \N__16456\,
            DOUT => \N__16455\,
            PACKAGEPIN => \SCLK1_wire\
        );

    \SCLK1_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__16457\,
            PADOUT => \N__16456\,
            PADIN => \N__16455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8992\,
            DIN0 => OPEN,
            DOUT0 => \N__14308\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCLK2_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__16448\,
            DIN => \N__16447\,
            DOUT => \N__16446\,
            PACKAGEPIN => \SCLK2_wire\
        );

    \SCLK2_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__16448\,
            PADOUT => \N__16447\,
            PADIN => \N__16446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8991\,
            DIN0 => OPEN,
            DOUT0 => \N__14307\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__16429\,
            I => \N__16426\
        );

    \I__3799\ : InMux
    port map (
            O => \N__16426\,
            I => \N__16423\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__16423\,
            I => \N__16420\
        );

    \I__3797\ : Span4Mux_h
    port map (
            O => \N__16420\,
            I => \N__16417\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__16417\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHGZ0\
        );

    \I__3795\ : InMux
    port map (
            O => \N__16414\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__3794\ : CascadeMux
    port map (
            O => \N__16411\,
            I => \N__16408\
        );

    \I__3793\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16404\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__16407\,
            I => \N__16398\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__16404\,
            I => \N__16391\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__16403\,
            I => \N__16388\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__16402\,
            I => \N__16385\
        );

    \I__3788\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16380\
        );

    \I__3787\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16377\
        );

    \I__3786\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16374\
        );

    \I__3785\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16371\
        );

    \I__3784\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16368\
        );

    \I__3783\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16365\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__16391\,
            I => \N__16361\
        );

    \I__3781\ : InMux
    port map (
            O => \N__16388\,
            I => \N__16356\
        );

    \I__3780\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16356\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__16384\,
            I => \N__16352\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__16383\,
            I => \N__16349\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__16380\,
            I => \N__16343\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__16377\,
            I => \N__16343\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__16374\,
            I => \N__16340\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__16371\,
            I => \N__16333\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__16368\,
            I => \N__16333\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__16365\,
            I => \N__16333\
        );

    \I__3771\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16330\
        );

    \I__3770\ : Sp12to4
    port map (
            O => \N__16361\,
            I => \N__16327\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__16356\,
            I => \N__16324\
        );

    \I__3768\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16319\
        );

    \I__3767\ : InMux
    port map (
            O => \N__16352\,
            I => \N__16319\
        );

    \I__3766\ : InMux
    port map (
            O => \N__16349\,
            I => \N__16316\
        );

    \I__3765\ : IoInMux
    port map (
            O => \N__16348\,
            I => \N__16313\
        );

    \I__3764\ : Span4Mux_v
    port map (
            O => \N__16343\,
            I => \N__16310\
        );

    \I__3763\ : Span4Mux_h
    port map (
            O => \N__16340\,
            I => \N__16303\
        );

    \I__3762\ : Span4Mux_v
    port map (
            O => \N__16333\,
            I => \N__16303\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__16330\,
            I => \N__16303\
        );

    \I__3760\ : Span12Mux_s10_h
    port map (
            O => \N__16327\,
            I => \N__16294\
        );

    \I__3759\ : Sp12to4
    port map (
            O => \N__16324\,
            I => \N__16294\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__16319\,
            I => \N__16294\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__16316\,
            I => \N__16294\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__16313\,
            I => \N__16291\
        );

    \I__3755\ : Span4Mux_h
    port map (
            O => \N__16310\,
            I => \N__16286\
        );

    \I__3754\ : Span4Mux_v
    port map (
            O => \N__16303\,
            I => \N__16286\
        );

    \I__3753\ : Span12Mux_v
    port map (
            O => \N__16294\,
            I => \N__16281\
        );

    \I__3752\ : Span12Mux_s1_v
    port map (
            O => \N__16291\,
            I => \N__16281\
        );

    \I__3751\ : Odrv4
    port map (
            O => \N__16286\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3750\ : Odrv12
    port map (
            O => \N__16281\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3749\ : CascadeMux
    port map (
            O => \N__16276\,
            I => \N__16273\
        );

    \I__3748\ : InMux
    port map (
            O => \N__16273\,
            I => \N__16270\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__16270\,
            I => \N__16267\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__16267\,
            I => \N__16264\
        );

    \I__3745\ : Odrv4
    port map (
            O => \N__16264\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6QZ0\
        );

    \I__3744\ : InMux
    port map (
            O => \N__16261\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__3743\ : InMux
    port map (
            O => \N__16258\,
            I => \N__16255\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__16255\,
            I => \N__16252\
        );

    \I__3741\ : Span4Mux_h
    port map (
            O => \N__16252\,
            I => \N__16249\
        );

    \I__3740\ : Odrv4
    port map (
            O => \N__16249\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8
        );

    \I__3739\ : InMux
    port map (
            O => \N__16246\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__3738\ : InMux
    port map (
            O => \N__16243\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7
        );

    \I__3737\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16237\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__16237\,
            I => \N__16232\
        );

    \I__3735\ : InMux
    port map (
            O => \N__16236\,
            I => \N__16229\
        );

    \I__3734\ : InMux
    port map (
            O => \N__16235\,
            I => \N__16226\
        );

    \I__3733\ : Span4Mux_v
    port map (
            O => \N__16232\,
            I => \N__16221\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__16229\,
            I => \N__16221\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__16226\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0\
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__16221\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0\
        );

    \I__3729\ : InMux
    port map (
            O => \N__16216\,
            I => \N__16213\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__16213\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\
        );

    \I__3727\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16204\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__16209\,
            I => \N__16195\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__16208\,
            I => \N__16192\
        );

    \I__3724\ : InMux
    port map (
            O => \N__16207\,
            I => \N__16187\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__16204\,
            I => \N__16180\
        );

    \I__3722\ : InMux
    port map (
            O => \N__16203\,
            I => \N__16173\
        );

    \I__3721\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16173\
        );

    \I__3720\ : InMux
    port map (
            O => \N__16201\,
            I => \N__16173\
        );

    \I__3719\ : InMux
    port map (
            O => \N__16200\,
            I => \N__16166\
        );

    \I__3718\ : InMux
    port map (
            O => \N__16199\,
            I => \N__16166\
        );

    \I__3717\ : InMux
    port map (
            O => \N__16198\,
            I => \N__16166\
        );

    \I__3716\ : InMux
    port map (
            O => \N__16195\,
            I => \N__16157\
        );

    \I__3715\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16157\
        );

    \I__3714\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16157\
        );

    \I__3713\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16157\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__16187\,
            I => \N__16148\
        );

    \I__3711\ : InMux
    port map (
            O => \N__16186\,
            I => \N__16139\
        );

    \I__3710\ : InMux
    port map (
            O => \N__16185\,
            I => \N__16139\
        );

    \I__3709\ : InMux
    port map (
            O => \N__16184\,
            I => \N__16139\
        );

    \I__3708\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16139\
        );

    \I__3707\ : Span4Mux_s2_h
    port map (
            O => \N__16180\,
            I => \N__16129\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__16173\,
            I => \N__16129\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__16166\,
            I => \N__16129\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16129\
        );

    \I__3703\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16126\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__16155\,
            I => \N__16123\
        );

    \I__3701\ : InMux
    port map (
            O => \N__16154\,
            I => \N__16120\
        );

    \I__3700\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16117\
        );

    \I__3699\ : InMux
    port map (
            O => \N__16152\,
            I => \N__16112\
        );

    \I__3698\ : InMux
    port map (
            O => \N__16151\,
            I => \N__16112\
        );

    \I__3697\ : Span4Mux_s3_h
    port map (
            O => \N__16148\,
            I => \N__16107\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__16139\,
            I => \N__16107\
        );

    \I__3695\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16104\
        );

    \I__3694\ : Span4Mux_h
    port map (
            O => \N__16129\,
            I => \N__16099\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__16126\,
            I => \N__16099\
        );

    \I__3692\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16096\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__16120\,
            I => \CO3_0\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__16117\,
            I => \CO3_0\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__16112\,
            I => \CO3_0\
        );

    \I__3688\ : Odrv4
    port map (
            O => \N__16107\,
            I => \CO3_0\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__16104\,
            I => \CO3_0\
        );

    \I__3686\ : Odrv4
    port map (
            O => \N__16099\,
            I => \CO3_0\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__16096\,
            I => \CO3_0\
        );

    \I__3684\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16078\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__16078\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i
        );

    \I__3682\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16063\
        );

    \I__3681\ : InMux
    port map (
            O => \N__16074\,
            I => \N__16063\
        );

    \I__3680\ : InMux
    port map (
            O => \N__16073\,
            I => \N__16063\
        );

    \I__3679\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16063\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__16063\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__3676\ : InMux
    port map (
            O => \N__16057\,
            I => \N__16054\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__16054\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKNZ0\
        );

    \I__3674\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16048\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__16048\,
            I => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\
        );

    \I__3672\ : InMux
    port map (
            O => \N__16045\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__3671\ : InMux
    port map (
            O => \N__16042\,
            I => \N__16039\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__16039\,
            I => \N__16036\
        );

    \I__3669\ : Odrv12
    port map (
            O => \N__16036\,
            I => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\
        );

    \I__3668\ : InMux
    port map (
            O => \N__16033\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__16030\,
            I => \N__16025\
        );

    \I__3666\ : InMux
    port map (
            O => \N__16029\,
            I => \N__15993\
        );

    \I__3665\ : InMux
    port map (
            O => \N__16028\,
            I => \N__15990\
        );

    \I__3664\ : InMux
    port map (
            O => \N__16025\,
            I => \N__15985\
        );

    \I__3663\ : InMux
    port map (
            O => \N__16024\,
            I => \N__15985\
        );

    \I__3662\ : InMux
    port map (
            O => \N__16023\,
            I => \N__15975\
        );

    \I__3661\ : InMux
    port map (
            O => \N__16022\,
            I => \N__15975\
        );

    \I__3660\ : InMux
    port map (
            O => \N__16021\,
            I => \N__15975\
        );

    \I__3659\ : InMux
    port map (
            O => \N__16020\,
            I => \N__15972\
        );

    \I__3658\ : InMux
    port map (
            O => \N__16019\,
            I => \N__15965\
        );

    \I__3657\ : InMux
    port map (
            O => \N__16018\,
            I => \N__15965\
        );

    \I__3656\ : InMux
    port map (
            O => \N__16017\,
            I => \N__15965\
        );

    \I__3655\ : InMux
    port map (
            O => \N__16016\,
            I => \N__15962\
        );

    \I__3654\ : InMux
    port map (
            O => \N__16015\,
            I => \N__15955\
        );

    \I__3653\ : InMux
    port map (
            O => \N__16014\,
            I => \N__15955\
        );

    \I__3652\ : InMux
    port map (
            O => \N__16013\,
            I => \N__15955\
        );

    \I__3651\ : InMux
    port map (
            O => \N__16012\,
            I => \N__15950\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16011\,
            I => \N__15950\
        );

    \I__3649\ : InMux
    port map (
            O => \N__16010\,
            I => \N__15945\
        );

    \I__3648\ : InMux
    port map (
            O => \N__16009\,
            I => \N__15945\
        );

    \I__3647\ : InMux
    port map (
            O => \N__16008\,
            I => \N__15936\
        );

    \I__3646\ : InMux
    port map (
            O => \N__16007\,
            I => \N__15936\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16006\,
            I => \N__15936\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16005\,
            I => \N__15936\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16004\,
            I => \N__15927\
        );

    \I__3642\ : InMux
    port map (
            O => \N__16003\,
            I => \N__15927\
        );

    \I__3641\ : InMux
    port map (
            O => \N__16002\,
            I => \N__15927\
        );

    \I__3640\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15927\
        );

    \I__3639\ : InMux
    port map (
            O => \N__16000\,
            I => \N__15920\
        );

    \I__3638\ : InMux
    port map (
            O => \N__15999\,
            I => \N__15920\
        );

    \I__3637\ : InMux
    port map (
            O => \N__15998\,
            I => \N__15920\
        );

    \I__3636\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15912\
        );

    \I__3635\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15912\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15905\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__15990\,
            I => \N__15905\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__15985\,
            I => \N__15905\
        );

    \I__3631\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15898\
        );

    \I__3630\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15898\
        );

    \I__3629\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15898\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__15975\,
            I => \N__15891\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__15972\,
            I => \N__15891\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__15965\,
            I => \N__15891\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__15962\,
            I => \N__15888\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__15955\,
            I => \N__15875\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__15950\,
            I => \N__15875\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__15945\,
            I => \N__15875\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__15936\,
            I => \N__15875\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__15927\,
            I => \N__15875\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__15920\,
            I => \N__15875\
        );

    \I__3618\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15870\
        );

    \I__3617\ : InMux
    port map (
            O => \N__15918\,
            I => \N__15870\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__15917\,
            I => \N__15863\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__15912\,
            I => \N__15854\
        );

    \I__3614\ : Span4Mux_h
    port map (
            O => \N__15905\,
            I => \N__15854\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__15898\,
            I => \N__15854\
        );

    \I__3612\ : Span4Mux_v
    port map (
            O => \N__15891\,
            I => \N__15851\
        );

    \I__3611\ : Span4Mux_h
    port map (
            O => \N__15888\,
            I => \N__15844\
        );

    \I__3610\ : Span4Mux_v
    port map (
            O => \N__15875\,
            I => \N__15844\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__15870\,
            I => \N__15844\
        );

    \I__3608\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15841\
        );

    \I__3607\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15828\
        );

    \I__3606\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15828\
        );

    \I__3605\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15828\
        );

    \I__3604\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15828\
        );

    \I__3603\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15828\
        );

    \I__3602\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15828\
        );

    \I__3601\ : Odrv4
    port map (
            O => \N__15854\,
            I => un5_rowlto1
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__15851\,
            I => un5_rowlto1
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__15844\,
            I => un5_rowlto1
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__15841\,
            I => un5_rowlto1
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__15828\,
            I => un5_rowlto1
        );

    \I__3596\ : CascadeMux
    port map (
            O => \N__15817\,
            I => \N__15809\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__15816\,
            I => \N__15800\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__15815\,
            I => \N__15797\
        );

    \I__3593\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15784\
        );

    \I__3592\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15784\
        );

    \I__3591\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15779\
        );

    \I__3590\ : InMux
    port map (
            O => \N__15809\,
            I => \N__15779\
        );

    \I__3589\ : InMux
    port map (
            O => \N__15808\,
            I => \N__15776\
        );

    \I__3588\ : InMux
    port map (
            O => \N__15807\,
            I => \N__15771\
        );

    \I__3587\ : InMux
    port map (
            O => \N__15806\,
            I => \N__15771\
        );

    \I__3586\ : InMux
    port map (
            O => \N__15805\,
            I => \N__15762\
        );

    \I__3585\ : InMux
    port map (
            O => \N__15804\,
            I => \N__15762\
        );

    \I__3584\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15762\
        );

    \I__3583\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15748\
        );

    \I__3582\ : InMux
    port map (
            O => \N__15797\,
            I => \N__15748\
        );

    \I__3581\ : InMux
    port map (
            O => \N__15796\,
            I => \N__15737\
        );

    \I__3580\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15737\
        );

    \I__3579\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15737\
        );

    \I__3578\ : InMux
    port map (
            O => \N__15793\,
            I => \N__15737\
        );

    \I__3577\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15737\
        );

    \I__3576\ : InMux
    port map (
            O => \N__15791\,
            I => \N__15734\
        );

    \I__3575\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15729\
        );

    \I__3574\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15729\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__15784\,
            I => \N__15723\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__15779\,
            I => \N__15723\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__15776\,
            I => \N__15718\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__15771\,
            I => \N__15718\
        );

    \I__3569\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15713\
        );

    \I__3568\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15713\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__15762\,
            I => \N__15710\
        );

    \I__3566\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15697\
        );

    \I__3565\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15697\
        );

    \I__3564\ : InMux
    port map (
            O => \N__15759\,
            I => \N__15697\
        );

    \I__3563\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15697\
        );

    \I__3562\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15697\
        );

    \I__3561\ : InMux
    port map (
            O => \N__15756\,
            I => \N__15697\
        );

    \I__3560\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15685\
        );

    \I__3559\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15685\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15753\,
            I => \N__15685\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__15748\,
            I => \N__15677\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__15737\,
            I => \N__15677\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__15734\,
            I => \N__15677\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__15729\,
            I => \N__15674\
        );

    \I__3553\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15671\
        );

    \I__3552\ : Span4Mux_v
    port map (
            O => \N__15723\,
            I => \N__15664\
        );

    \I__3551\ : Span4Mux_v
    port map (
            O => \N__15718\,
            I => \N__15664\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__15713\,
            I => \N__15664\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__15710\,
            I => \N__15659\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__15697\,
            I => \N__15659\
        );

    \I__3547\ : InMux
    port map (
            O => \N__15696\,
            I => \N__15648\
        );

    \I__3546\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15648\
        );

    \I__3545\ : InMux
    port map (
            O => \N__15694\,
            I => \N__15648\
        );

    \I__3544\ : InMux
    port map (
            O => \N__15693\,
            I => \N__15648\
        );

    \I__3543\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15648\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__15685\,
            I => \N__15645\
        );

    \I__3541\ : InMux
    port map (
            O => \N__15684\,
            I => \N__15642\
        );

    \I__3540\ : Span4Mux_h
    port map (
            O => \N__15677\,
            I => \N__15639\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__15674\,
            I => un5_rowlto0
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__15671\,
            I => un5_rowlto0
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__15664\,
            I => un5_rowlto0
        );

    \I__3536\ : Odrv4
    port map (
            O => \N__15659\,
            I => un5_rowlto0
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__15648\,
            I => un5_rowlto0
        );

    \I__3534\ : Odrv12
    port map (
            O => \N__15645\,
            I => un5_rowlto0
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__15642\,
            I => un5_rowlto0
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__15639\,
            I => un5_rowlto0
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__15622\,
            I => \un5_rowlto1_cascade_\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__15618\,
            I => \N__15610\
        );

    \I__3528\ : InMux
    port map (
            O => \N__15617\,
            I => \N__15605\
        );

    \I__3527\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15602\
        );

    \I__3526\ : InMux
    port map (
            O => \N__15613\,
            I => \N__15595\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15595\
        );

    \I__3524\ : InMux
    port map (
            O => \N__15609\,
            I => \N__15595\
        );

    \I__3523\ : InMux
    port map (
            O => \N__15608\,
            I => \N__15581\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__15605\,
            I => \N__15574\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__15602\,
            I => \N__15571\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15568\
        );

    \I__3519\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15563\
        );

    \I__3518\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15563\
        );

    \I__3517\ : InMux
    port map (
            O => \N__15592\,
            I => \N__15560\
        );

    \I__3516\ : InMux
    port map (
            O => \N__15591\,
            I => \N__15555\
        );

    \I__3515\ : InMux
    port map (
            O => \N__15590\,
            I => \N__15555\
        );

    \I__3514\ : InMux
    port map (
            O => \N__15589\,
            I => \N__15552\
        );

    \I__3513\ : InMux
    port map (
            O => \N__15588\,
            I => \N__15549\
        );

    \I__3512\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15546\
        );

    \I__3511\ : InMux
    port map (
            O => \N__15586\,
            I => \N__15541\
        );

    \I__3510\ : InMux
    port map (
            O => \N__15585\,
            I => \N__15538\
        );

    \I__3509\ : InMux
    port map (
            O => \N__15584\,
            I => \N__15535\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__15581\,
            I => \N__15532\
        );

    \I__3507\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15529\
        );

    \I__3506\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15526\
        );

    \I__3505\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15521\
        );

    \I__3504\ : InMux
    port map (
            O => \N__15577\,
            I => \N__15521\
        );

    \I__3503\ : Span4Mux_s1_h
    port map (
            O => \N__15574\,
            I => \N__15512\
        );

    \I__3502\ : Span4Mux_v
    port map (
            O => \N__15571\,
            I => \N__15512\
        );

    \I__3501\ : Span4Mux_v
    port map (
            O => \N__15568\,
            I => \N__15512\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__15563\,
            I => \N__15512\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__15560\,
            I => \N__15505\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__15555\,
            I => \N__15505\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__15552\,
            I => \N__15505\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__15549\,
            I => \N__15500\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__15546\,
            I => \N__15500\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__15545\,
            I => \N__15496\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__15544\,
            I => \N__15493\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15489\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__15538\,
            I => \N__15486\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15535\,
            I => \N__15475\
        );

    \I__3489\ : Span4Mux_h
    port map (
            O => \N__15532\,
            I => \N__15475\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__15529\,
            I => \N__15475\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__15526\,
            I => \N__15475\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__15521\,
            I => \N__15475\
        );

    \I__3485\ : Span4Mux_h
    port map (
            O => \N__15512\,
            I => \N__15472\
        );

    \I__3484\ : Span4Mux_v
    port map (
            O => \N__15505\,
            I => \N__15467\
        );

    \I__3483\ : Span4Mux_h
    port map (
            O => \N__15500\,
            I => \N__15467\
        );

    \I__3482\ : InMux
    port map (
            O => \N__15499\,
            I => \N__15464\
        );

    \I__3481\ : InMux
    port map (
            O => \N__15496\,
            I => \N__15457\
        );

    \I__3480\ : InMux
    port map (
            O => \N__15493\,
            I => \N__15457\
        );

    \I__3479\ : InMux
    port map (
            O => \N__15492\,
            I => \N__15457\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__15489\,
            I => un5_rowlto3
        );

    \I__3477\ : Odrv12
    port map (
            O => \N__15486\,
            I => un5_rowlto3
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__15475\,
            I => un5_rowlto3
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__15472\,
            I => un5_rowlto3
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__15467\,
            I => un5_rowlto3
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__15464\,
            I => un5_rowlto3
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__15457\,
            I => un5_rowlto3
        );

    \I__3471\ : InMux
    port map (
            O => \N__15442\,
            I => \N__15439\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__15439\,
            I => \N__15436\
        );

    \I__3469\ : Span4Mux_h
    port map (
            O => \N__15436\,
            I => \N__15433\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__15433\,
            I => un116_pixel_2_am_0
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__15430\,
            I => \N__15426\
        );

    \I__3466\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15421\
        );

    \I__3465\ : InMux
    port map (
            O => \N__15426\,
            I => \N__15421\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__15421\,
            I => \N__15418\
        );

    \I__3463\ : Span4Mux_s1_h
    port map (
            O => \N__15418\,
            I => \N__15415\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__15415\,
            I => if_generate_plus_mult1_un68_sum_cry_3_s
        );

    \I__3461\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15409\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__15409\,
            I => if_generate_plus_mult1_un75_sum_axb_4_l_fx
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__15406\,
            I => \N__15390\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__15405\,
            I => \N__15386\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__15404\,
            I => \N__15377\
        );

    \I__3456\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15368\
        );

    \I__3455\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15368\
        );

    \I__3454\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15368\
        );

    \I__3453\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15357\
        );

    \I__3452\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15357\
        );

    \I__3451\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15357\
        );

    \I__3450\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15357\
        );

    \I__3449\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15357\
        );

    \I__3448\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15349\
        );

    \I__3447\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15349\
        );

    \I__3446\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15338\
        );

    \I__3445\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15338\
        );

    \I__3444\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15338\
        );

    \I__3443\ : InMux
    port map (
            O => \N__15386\,
            I => \N__15338\
        );

    \I__3442\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15338\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__15384\,
            I => \N__15330\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__15383\,
            I => \N__15327\
        );

    \I__3439\ : InMux
    port map (
            O => \N__15382\,
            I => \N__15323\
        );

    \I__3438\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15312\
        );

    \I__3437\ : InMux
    port map (
            O => \N__15380\,
            I => \N__15312\
        );

    \I__3436\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15312\
        );

    \I__3435\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15312\
        );

    \I__3434\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15312\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__15368\,
            I => \N__15309\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__15357\,
            I => \N__15306\
        );

    \I__3431\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15303\
        );

    \I__3430\ : InMux
    port map (
            O => \N__15355\,
            I => \N__15289\
        );

    \I__3429\ : InMux
    port map (
            O => \N__15354\,
            I => \N__15289\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__15349\,
            I => \N__15282\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__15338\,
            I => \N__15282\
        );

    \I__3426\ : InMux
    port map (
            O => \N__15337\,
            I => \N__15277\
        );

    \I__3425\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15277\
        );

    \I__3424\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15272\
        );

    \I__3423\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15272\
        );

    \I__3422\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15269\
        );

    \I__3421\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15262\
        );

    \I__3420\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15262\
        );

    \I__3419\ : InMux
    port map (
            O => \N__15326\,
            I => \N__15262\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__15323\,
            I => \N__15259\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__15312\,
            I => \N__15250\
        );

    \I__3416\ : Span4Mux_v
    port map (
            O => \N__15309\,
            I => \N__15250\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__15306\,
            I => \N__15250\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15250\
        );

    \I__3413\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15244\
        );

    \I__3412\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15244\
        );

    \I__3411\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15241\
        );

    \I__3410\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15234\
        );

    \I__3409\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15234\
        );

    \I__3408\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15234\
        );

    \I__3407\ : InMux
    port map (
            O => \N__15296\,
            I => \N__15229\
        );

    \I__3406\ : InMux
    port map (
            O => \N__15295\,
            I => \N__15229\
        );

    \I__3405\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15226\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__15289\,
            I => \N__15223\
        );

    \I__3403\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15220\
        );

    \I__3402\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15217\
        );

    \I__3401\ : Span4Mux_v
    port map (
            O => \N__15282\,
            I => \N__15214\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__15277\,
            I => \N__15205\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__15272\,
            I => \N__15205\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__15269\,
            I => \N__15205\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__15262\,
            I => \N__15205\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__15259\,
            I => \N__15200\
        );

    \I__3395\ : Span4Mux_h
    port map (
            O => \N__15250\,
            I => \N__15200\
        );

    \I__3394\ : InMux
    port map (
            O => \N__15249\,
            I => \N__15197\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__15244\,
            I => \N__15190\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__15241\,
            I => \N__15190\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__15234\,
            I => \N__15190\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__15229\,
            I => un5_rowlto2
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__15226\,
            I => un5_rowlto2
        );

    \I__3388\ : Odrv12
    port map (
            O => \N__15223\,
            I => un5_rowlto2
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__15220\,
            I => un5_rowlto2
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__15217\,
            I => un5_rowlto2
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__15214\,
            I => un5_rowlto2
        );

    \I__3384\ : Odrv4
    port map (
            O => \N__15205\,
            I => un5_rowlto2
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__15200\,
            I => un5_rowlto2
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__15197\,
            I => un5_rowlto2
        );

    \I__3381\ : Odrv12
    port map (
            O => \N__15190\,
            I => un5_rowlto2
        );

    \I__3380\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15166\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__15166\,
            I => un5_rowlto2_i
        );

    \I__3378\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15159\
        );

    \I__3377\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15156\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__15159\,
            I => \N__15152\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__15156\,
            I => \N__15149\
        );

    \I__3374\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15145\
        );

    \I__3373\ : Span4Mux_v
    port map (
            O => \N__15152\,
            I => \N__15140\
        );

    \I__3372\ : Span4Mux_s1_h
    port map (
            O => \N__15149\,
            I => \N__15140\
        );

    \I__3371\ : InMux
    port map (
            O => \N__15148\,
            I => \N__15137\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__15145\,
            I => \N__15134\
        );

    \I__3369\ : Span4Mux_h
    port map (
            O => \N__15140\,
            I => \N__15131\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__15137\,
            I => \N__15126\
        );

    \I__3367\ : Span4Mux_v
    port map (
            O => \N__15134\,
            I => \N__15126\
        );

    \I__3366\ : Odrv4
    port map (
            O => \N__15131\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__3365\ : Odrv4
    port map (
            O => \N__15126\,
            I => charx_if_generate_plus_mult1_un68_sum
        );

    \I__3364\ : CascadeMux
    port map (
            O => \N__15121\,
            I => \N__15118\
        );

    \I__3363\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15115\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__15115\,
            I => \N__15112\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__15112\,
            I => \column_1_if_generate_plus_mult1_un75_sum_iZ0\
        );

    \I__3360\ : InMux
    port map (
            O => \N__15109\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__15106\,
            I => \N__15103\
        );

    \I__3358\ : InMux
    port map (
            O => \N__15103\,
            I => \N__15099\
        );

    \I__3357\ : InMux
    port map (
            O => \N__15102\,
            I => \N__15094\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__15099\,
            I => \N__15090\
        );

    \I__3355\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15085\
        );

    \I__3354\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15085\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__15094\,
            I => \N__15082\
        );

    \I__3352\ : CascadeMux
    port map (
            O => \N__15093\,
            I => \N__15078\
        );

    \I__3351\ : Span4Mux_v
    port map (
            O => \N__15090\,
            I => \N__15072\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__15085\,
            I => \N__15072\
        );

    \I__3349\ : Span4Mux_s1_h
    port map (
            O => \N__15082\,
            I => \N__15069\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15066\
        );

    \I__3347\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15062\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15077\,
            I => \N__15059\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__15072\,
            I => \N__15056\
        );

    \I__3344\ : Span4Mux_h
    port map (
            O => \N__15069\,
            I => \N__15051\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__15066\,
            I => \N__15051\
        );

    \I__3342\ : InMux
    port map (
            O => \N__15065\,
            I => \N__15048\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__15062\,
            I => \N__15045\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__15059\,
            I => charx_if_generate_plus_mult1_un26_sum
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__15056\,
            I => charx_if_generate_plus_mult1_un26_sum
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__15051\,
            I => charx_if_generate_plus_mult1_un26_sum
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__15048\,
            I => charx_if_generate_plus_mult1_un26_sum
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__15045\,
            I => charx_if_generate_plus_mult1_un26_sum
        );

    \I__3335\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15031\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__15031\,
            I => \G_346\
        );

    \I__3333\ : InMux
    port map (
            O => \N__15028\,
            I => column_1_if_generate_plus_mult1_un82_sum_cry_4
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__15025\,
            I => \un5_rowlto0_cascade_\
        );

    \I__3331\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15019\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__15019\,
            I => \un116_pixel_1_bmZ0Z_1\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__15016\,
            I => \N__15004\
        );

    \I__3328\ : CascadeMux
    port map (
            O => \N__15015\,
            I => \N__15000\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__15014\,
            I => \N__14996\
        );

    \I__3326\ : InMux
    port map (
            O => \N__15013\,
            I => \N__14991\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__15012\,
            I => \N__14988\
        );

    \I__3324\ : InMux
    port map (
            O => \N__15011\,
            I => \N__14977\
        );

    \I__3323\ : InMux
    port map (
            O => \N__15010\,
            I => \N__14977\
        );

    \I__3322\ : InMux
    port map (
            O => \N__15009\,
            I => \N__14977\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__15008\,
            I => \N__14971\
        );

    \I__3320\ : InMux
    port map (
            O => \N__15007\,
            I => \N__14968\
        );

    \I__3319\ : InMux
    port map (
            O => \N__15004\,
            I => \N__14965\
        );

    \I__3318\ : InMux
    port map (
            O => \N__15003\,
            I => \N__14960\
        );

    \I__3317\ : InMux
    port map (
            O => \N__15000\,
            I => \N__14960\
        );

    \I__3316\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14955\
        );

    \I__3315\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14955\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__14995\,
            I => \N__14951\
        );

    \I__3313\ : InMux
    port map (
            O => \N__14994\,
            I => \N__14946\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__14991\,
            I => \N__14943\
        );

    \I__3311\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14940\
        );

    \I__3310\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14935\
        );

    \I__3309\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14935\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14985\,
            I => \N__14930\
        );

    \I__3307\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14930\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__14977\,
            I => \N__14927\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__14976\,
            I => \N__14924\
        );

    \I__3304\ : CascadeMux
    port map (
            O => \N__14975\,
            I => \N__14921\
        );

    \I__3303\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14917\
        );

    \I__3302\ : InMux
    port map (
            O => \N__14971\,
            I => \N__14914\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__14968\,
            I => \N__14909\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__14965\,
            I => \N__14909\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__14960\,
            I => \N__14904\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__14955\,
            I => \N__14904\
        );

    \I__3297\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14897\
        );

    \I__3296\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14894\
        );

    \I__3295\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14889\
        );

    \I__3294\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14889\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__14946\,
            I => \N__14886\
        );

    \I__3292\ : Span4Mux_s2_h
    port map (
            O => \N__14943\,
            I => \N__14883\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__14940\,
            I => \N__14874\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__14935\,
            I => \N__14874\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__14930\,
            I => \N__14874\
        );

    \I__3288\ : Span4Mux_s1_h
    port map (
            O => \N__14927\,
            I => \N__14874\
        );

    \I__3287\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14871\
        );

    \I__3286\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14868\
        );

    \I__3285\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14865\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__14917\,
            I => \N__14862\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__14914\,
            I => \N__14859\
        );

    \I__3282\ : Span4Mux_h
    port map (
            O => \N__14909\,
            I => \N__14856\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__14904\,
            I => \N__14853\
        );

    \I__3280\ : InMux
    port map (
            O => \N__14903\,
            I => \N__14850\
        );

    \I__3279\ : InMux
    port map (
            O => \N__14902\,
            I => \N__14843\
        );

    \I__3278\ : InMux
    port map (
            O => \N__14901\,
            I => \N__14843\
        );

    \I__3277\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14843\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__14897\,
            I => \N__14836\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__14894\,
            I => \N__14836\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__14889\,
            I => \N__14836\
        );

    \I__3273\ : Span4Mux_h
    port map (
            O => \N__14886\,
            I => \N__14829\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__14883\,
            I => \N__14829\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__14874\,
            I => \N__14829\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__14871\,
            I => \N__14822\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__14868\,
            I => \N__14822\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__14865\,
            I => \N__14822\
        );

    \I__3267\ : Odrv4
    port map (
            O => \N__14862\,
            I => \beamYZ0Z_1\
        );

    \I__3266\ : Odrv12
    port map (
            O => \N__14859\,
            I => \beamYZ0Z_1\
        );

    \I__3265\ : Odrv4
    port map (
            O => \N__14856\,
            I => \beamYZ0Z_1\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__14853\,
            I => \beamYZ0Z_1\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__14850\,
            I => \beamYZ0Z_1\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__14843\,
            I => \beamYZ0Z_1\
        );

    \I__3261\ : Odrv12
    port map (
            O => \N__14836\,
            I => \beamYZ0Z_1\
        );

    \I__3260\ : Odrv4
    port map (
            O => \N__14829\,
            I => \beamYZ0Z_1\
        );

    \I__3259\ : Odrv12
    port map (
            O => \N__14822\,
            I => \beamYZ0Z_1\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__14803\,
            I => \un116_pixel_1_bmZ0Z_1_cascade_\
        );

    \I__3257\ : InMux
    port map (
            O => \N__14800\,
            I => \N__14797\
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__14797\,
            I => \N__14794\
        );

    \I__3255\ : Span4Mux_h
    port map (
            O => \N__14794\,
            I => \N__14791\
        );

    \I__3254\ : Odrv4
    port map (
            O => \N__14791\,
            I => \beamY_RNIV622TRZ0Z_1\
        );

    \I__3253\ : InMux
    port map (
            O => \N__14788\,
            I => \N__14785\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__14785\,
            I => \N__14782\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__14782\,
            I => un116_pixel_2_ns_1_4
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__14779\,
            I => \N__14770\
        );

    \I__3249\ : CascadeMux
    port map (
            O => \N__14778\,
            I => \N__14762\
        );

    \I__3248\ : CascadeMux
    port map (
            O => \N__14777\,
            I => \N__14754\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__14776\,
            I => \N__14747\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__14775\,
            I => \N__14738\
        );

    \I__3245\ : CascadeMux
    port map (
            O => \N__14774\,
            I => \N__14733\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__14773\,
            I => \N__14730\
        );

    \I__3243\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14726\
        );

    \I__3242\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14723\
        );

    \I__3241\ : InMux
    port map (
            O => \N__14768\,
            I => \N__14714\
        );

    \I__3240\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14714\
        );

    \I__3239\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14714\
        );

    \I__3238\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14714\
        );

    \I__3237\ : InMux
    port map (
            O => \N__14762\,
            I => \N__14709\
        );

    \I__3236\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14709\
        );

    \I__3235\ : InMux
    port map (
            O => \N__14760\,
            I => \N__14706\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__14759\,
            I => \N__14703\
        );

    \I__3233\ : InMux
    port map (
            O => \N__14758\,
            I => \N__14695\
        );

    \I__3232\ : InMux
    port map (
            O => \N__14757\,
            I => \N__14695\
        );

    \I__3231\ : InMux
    port map (
            O => \N__14754\,
            I => \N__14695\
        );

    \I__3230\ : InMux
    port map (
            O => \N__14753\,
            I => \N__14690\
        );

    \I__3229\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14690\
        );

    \I__3228\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14687\
        );

    \I__3227\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14684\
        );

    \I__3226\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14681\
        );

    \I__3225\ : InMux
    port map (
            O => \N__14746\,
            I => \N__14676\
        );

    \I__3224\ : InMux
    port map (
            O => \N__14745\,
            I => \N__14676\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__14744\,
            I => \N__14673\
        );

    \I__3222\ : InMux
    port map (
            O => \N__14743\,
            I => \N__14666\
        );

    \I__3221\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14666\
        );

    \I__3220\ : InMux
    port map (
            O => \N__14741\,
            I => \N__14666\
        );

    \I__3219\ : InMux
    port map (
            O => \N__14738\,
            I => \N__14657\
        );

    \I__3218\ : InMux
    port map (
            O => \N__14737\,
            I => \N__14657\
        );

    \I__3217\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14657\
        );

    \I__3216\ : InMux
    port map (
            O => \N__14733\,
            I => \N__14657\
        );

    \I__3215\ : InMux
    port map (
            O => \N__14730\,
            I => \N__14652\
        );

    \I__3214\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14652\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14645\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__14723\,
            I => \N__14645\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__14714\,
            I => \N__14645\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__14709\,
            I => \N__14642\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__14706\,
            I => \N__14638\
        );

    \I__3208\ : InMux
    port map (
            O => \N__14703\,
            I => \N__14635\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__14702\,
            I => \N__14631\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__14695\,
            I => \N__14627\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__14690\,
            I => \N__14622\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__14687\,
            I => \N__14622\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14617\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__14681\,
            I => \N__14617\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__14676\,
            I => \N__14614\
        );

    \I__3200\ : InMux
    port map (
            O => \N__14673\,
            I => \N__14611\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__14666\,
            I => \N__14608\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__14657\,
            I => \N__14599\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__14652\,
            I => \N__14599\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__14645\,
            I => \N__14599\
        );

    \I__3195\ : Span4Mux_s1_h
    port map (
            O => \N__14642\,
            I => \N__14599\
        );

    \I__3194\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14596\
        );

    \I__3193\ : Span12Mux_s5_h
    port map (
            O => \N__14638\,
            I => \N__14593\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__14635\,
            I => \N__14590\
        );

    \I__3191\ : InMux
    port map (
            O => \N__14634\,
            I => \N__14587\
        );

    \I__3190\ : InMux
    port map (
            O => \N__14631\,
            I => \N__14582\
        );

    \I__3189\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14582\
        );

    \I__3188\ : Span4Mux_h
    port map (
            O => \N__14627\,
            I => \N__14577\
        );

    \I__3187\ : Span4Mux_h
    port map (
            O => \N__14622\,
            I => \N__14577\
        );

    \I__3186\ : Span4Mux_h
    port map (
            O => \N__14617\,
            I => \N__14574\
        );

    \I__3185\ : Span4Mux_v
    port map (
            O => \N__14614\,
            I => \N__14569\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__14611\,
            I => \N__14569\
        );

    \I__3183\ : Span4Mux_v
    port map (
            O => \N__14608\,
            I => \N__14564\
        );

    \I__3182\ : Span4Mux_h
    port map (
            O => \N__14599\,
            I => \N__14564\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__14596\,
            I => \beamYZ0Z_0\
        );

    \I__3180\ : Odrv12
    port map (
            O => \N__14593\,
            I => \beamYZ0Z_0\
        );

    \I__3179\ : Odrv4
    port map (
            O => \N__14590\,
            I => \beamYZ0Z_0\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__14587\,
            I => \beamYZ0Z_0\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__14582\,
            I => \beamYZ0Z_0\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__14577\,
            I => \beamYZ0Z_0\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__14574\,
            I => \beamYZ0Z_0\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__14569\,
            I => \beamYZ0Z_0\
        );

    \I__3173\ : Odrv4
    port map (
            O => \N__14564\,
            I => \beamYZ0Z_0\
        );

    \I__3172\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__14542\,
            I => \N__14539\
        );

    \I__3170\ : Odrv4
    port map (
            O => \N__14539\,
            I => \beamY_RNIITCG3J3Z0Z_0\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__14536\,
            I => \N__14533\
        );

    \I__3168\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14530\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__14530\,
            I => \N__14527\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__14527\,
            I => \column_1_if_generate_plus_mult1_un68_sum_iZ0\
        );

    \I__3165\ : InMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__14521\,
            I => if_generate_plus_mult1_un75_sum_cry_2_s
        );

    \I__3163\ : InMux
    port map (
            O => \N__14518\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__14515\,
            I => \N__14512\
        );

    \I__3161\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14509\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__14509\,
            I => \N__14506\
        );

    \I__3159\ : Odrv12
    port map (
            O => \N__14506\,
            I => if_generate_plus_mult1_un68_sum_cry_2_s
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__14503\,
            I => \N__14500\
        );

    \I__3157\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14497\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__14497\,
            I => if_generate_plus_mult1_un75_sum_cry_3_s
        );

    \I__3155\ : InMux
    port map (
            O => \N__14494\,
            I => column_1_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__3154\ : InMux
    port map (
            O => \N__14491\,
            I => \N__14488\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__14488\,
            I => \un116_pixel_2_bmZ0Z_5\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__14485\,
            I => \un114_pixel_7_1_7__N_9_cascade_\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__14482\,
            I => \un114_pixel_1_0_3__un116_pixel_3_ns_1Z0Z_0_cascade_\
        );

    \I__3150\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14476\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__14476\,
            I => \un114_pixel_6_1_5__N_8\
        );

    \I__3148\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14470\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__14470\,
            I => \N__14467\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__14467\,
            I => \N__14464\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__14464\,
            I => \N_371\
        );

    \I__3144\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14458\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__14458\,
            I => \N__14455\
        );

    \I__3142\ : Odrv4
    port map (
            O => \N__14455\,
            I => \beamY_RNIJUCG3J3Z0Z_1\
        );

    \I__3141\ : InMux
    port map (
            O => \N__14452\,
            I => \N__14447\
        );

    \I__3140\ : InMux
    port map (
            O => \N__14451\,
            I => \N__14441\
        );

    \I__3139\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14438\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__14447\,
            I => \N__14435\
        );

    \I__3137\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14430\
        );

    \I__3136\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14430\
        );

    \I__3135\ : InMux
    port map (
            O => \N__14444\,
            I => \N__14427\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__14441\,
            I => \N__14420\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__14438\,
            I => \N__14420\
        );

    \I__3132\ : Span4Mux_s3_h
    port map (
            O => \N__14435\,
            I => \N__14415\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__14430\,
            I => \N__14415\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__14427\,
            I => \N__14412\
        );

    \I__3129\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14407\
        );

    \I__3128\ : InMux
    port map (
            O => \N__14425\,
            I => \N__14407\
        );

    \I__3127\ : Span4Mux_v
    port map (
            O => \N__14420\,
            I => \N__14398\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__14415\,
            I => \N__14398\
        );

    \I__3125\ : Span4Mux_s3_h
    port map (
            O => \N__14412\,
            I => \N__14398\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__14407\,
            I => \N__14398\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__14398\,
            I => charx_if_generate_plus_mult1_un75_sum
        );

    \I__3122\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14392\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__14392\,
            I => \G_345\
        );

    \I__3120\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__3119\ : InMux
    port map (
            O => \N__14388\,
            I => \N__14383\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__14383\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8
        );

    \I__3117\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14377\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__14377\,
            I => \N__14374\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__14374\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8
        );

    \I__3114\ : InMux
    port map (
            O => \N__14371\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__3113\ : InMux
    port map (
            O => \N__14368\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7
        );

    \I__3112\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14362\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__14362\,
            I => \N__14357\
        );

    \I__3110\ : InMux
    port map (
            O => \N__14361\,
            I => \N__14354\
        );

    \I__3109\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14351\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__14357\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__14354\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__14351\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__14344\,
            I => \N__14341\
        );

    \I__3104\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14338\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__14338\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i
        );

    \I__3102\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14332\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__14332\,
            I => \N__14329\
        );

    \I__3100\ : Glb2LocalMux
    port map (
            O => \N__14329\,
            I => \N__14314\
        );

    \I__3099\ : ClkMux
    port map (
            O => \N__14328\,
            I => \N__14314\
        );

    \I__3098\ : ClkMux
    port map (
            O => \N__14327\,
            I => \N__14314\
        );

    \I__3097\ : ClkMux
    port map (
            O => \N__14326\,
            I => \N__14314\
        );

    \I__3096\ : ClkMux
    port map (
            O => \N__14325\,
            I => \N__14314\
        );

    \I__3095\ : GlobalMux
    port map (
            O => \N__14314\,
            I => \N__14311\
        );

    \I__3094\ : gio2CtrlBuf
    port map (
            O => \N__14311\,
            I => \Clock12MHz_c_g\
        );

    \I__3093\ : IoInMux
    port map (
            O => \N__14308\,
            I => \N__14303\
        );

    \I__3092\ : IoInMux
    port map (
            O => \N__14307\,
            I => \N__14300\
        );

    \I__3091\ : IoInMux
    port map (
            O => \N__14306\,
            I => \N__14297\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__14303\,
            I => \N__14292\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__14300\,
            I => \N__14292\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__14297\,
            I => \N__14289\
        );

    \I__3087\ : Span12Mux_s11_v
    port map (
            O => \N__14292\,
            I => \N__14286\
        );

    \I__3086\ : Span12Mux_s10_h
    port map (
            O => \N__14289\,
            I => \N__14283\
        );

    \I__3085\ : Odrv12
    port map (
            O => \N__14286\,
            I => \GB_BUFFER_Clock12MHz_c_g_THRU_CO\
        );

    \I__3084\ : Odrv12
    port map (
            O => \N__14283\,
            I => \GB_BUFFER_Clock12MHz_c_g_THRU_CO\
        );

    \I__3083\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14275\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__14275\,
            I => \N__14272\
        );

    \I__3081\ : Odrv4
    port map (
            O => \N__14272\,
            I => \N_1557_0\
        );

    \I__3080\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14266\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__14266\,
            I => \N__14263\
        );

    \I__3078\ : Odrv12
    port map (
            O => \N__14263\,
            I => \N_41_0_0_0\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__14260\,
            I => \N__14257\
        );

    \I__3076\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14250\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__14256\,
            I => \N__14247\
        );

    \I__3074\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14241\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__14254\,
            I => \N__14234\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__14253\,
            I => \N__14231\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__14250\,
            I => \N__14228\
        );

    \I__3070\ : InMux
    port map (
            O => \N__14247\,
            I => \N__14225\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__14246\,
            I => \N__14222\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__14245\,
            I => \N__14218\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__14244\,
            I => \N__14214\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14211\
        );

    \I__3065\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14206\
        );

    \I__3064\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14206\
        );

    \I__3063\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14203\
        );

    \I__3062\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14196\
        );

    \I__3061\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14196\
        );

    \I__3060\ : InMux
    port map (
            O => \N__14231\,
            I => \N__14196\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__14228\,
            I => \N__14191\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__14225\,
            I => \N__14191\
        );

    \I__3057\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14184\
        );

    \I__3056\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14184\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14184\
        );

    \I__3054\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14179\
        );

    \I__3053\ : InMux
    port map (
            O => \N__14214\,
            I => \N__14179\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__14211\,
            I => \N_563\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N_563\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__14203\,
            I => \N_563\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__14196\,
            I => \N_563\
        );

    \I__3048\ : Odrv4
    port map (
            O => \N__14191\,
            I => \N_563\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__14184\,
            I => \N_563\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__14179\,
            I => \N_563\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__14164\,
            I => \un116_pixel_5_bmZ0Z_5_cascade_\
        );

    \I__3044\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14158\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__14155\,
            I => \N__14152\
        );

    \I__3041\ : Odrv4
    port map (
            O => \N__14152\,
            I => un116_pixel_6_ns_1_5
        );

    \I__3040\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14146\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__14146\,
            I => if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__14143\,
            I => \N__14140\
        );

    \I__3037\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14137\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__14137\,
            I => \N_858_i\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__14134\,
            I => \N__14131\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14131\,
            I => \N__14128\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__14128\,
            I => \N__14125\
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__14125\,
            I => column_1_if_generate_plus_mult1_un47_sum1_3
        );

    \I__3031\ : InMux
    port map (
            O => \N__14122\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_2
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__14119\,
            I => \N__14116\
        );

    \I__3029\ : InMux
    port map (
            O => \N__14116\,
            I => \N__14113\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__14113\,
            I => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx
        );

    \I__3027\ : InMux
    port map (
            O => \N__14110\,
            I => \N__14107\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__14107\,
            I => column_1_if_generate_plus_mult1_un47_sum1_4
        );

    \I__3025\ : InMux
    port map (
            O => \N__14104\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_3
        );

    \I__3024\ : InMux
    port map (
            O => \N__14101\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_4
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__14098\,
            I => \N__14094\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__14097\,
            I => \N__14090\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14086\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14093\,
            I => \N__14079\
        );

    \I__3019\ : InMux
    port map (
            O => \N__14090\,
            I => \N__14079\
        );

    \I__3018\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14079\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__14086\,
            I => column_1_if_generate_plus_mult1_un47_sum1_5
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__14079\,
            I => column_1_if_generate_plus_mult1_un47_sum1_5
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__14074\,
            I => \N__14070\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__14073\,
            I => \N__14067\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14070\,
            I => \N__14062\
        );

    \I__3012\ : InMux
    port map (
            O => \N__14067\,
            I => \N__14062\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__14062\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8
        );

    \I__3010\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14054\
        );

    \I__3009\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14049\
        );

    \I__3008\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14049\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__14054\,
            I => \N__14043\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__14049\,
            I => \N__14043\
        );

    \I__3005\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14040\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__14043\,
            I => \N__14033\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__14040\,
            I => \N__14033\
        );

    \I__3002\ : InMux
    port map (
            O => \N__14039\,
            I => \N__14025\
        );

    \I__3001\ : InMux
    port map (
            O => \N__14038\,
            I => \N__14025\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__14033\,
            I => \N__14022\
        );

    \I__2999\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14017\
        );

    \I__2998\ : InMux
    port map (
            O => \N__14031\,
            I => \N__14017\
        );

    \I__2997\ : InMux
    port map (
            O => \N__14030\,
            I => \N__14014\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__14025\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2995\ : Odrv4
    port map (
            O => \N__14022\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__14017\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__14014\,
            I => charx_if_generate_plus_mult1_un33_sum
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__14005\,
            I => \N__14000\
        );

    \I__2991\ : InMux
    port map (
            O => \N__14004\,
            I => \N__13995\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14003\,
            I => \N__13995\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13992\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__13995\,
            I => \N__13989\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__13992\,
            I => \N_66\
        );

    \I__2986\ : Odrv4
    port map (
            O => \N__13989\,
            I => \N_66\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__13984\,
            I => \N__13981\
        );

    \I__2984\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13978\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__13978\,
            I => \N__13975\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__13975\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5LZ0\
        );

    \I__2981\ : InMux
    port map (
            O => \N__13972\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2980\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13966\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__13966\,
            I => \N__13963\
        );

    \I__2978\ : Odrv4
    port map (
            O => \N__13963\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7JZ0Z31\
        );

    \I__2977\ : InMux
    port map (
            O => \N__13960\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__2976\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13954\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__13954\,
            I => \N__13951\
        );

    \I__2974\ : Odrv12
    port map (
            O => \N__13951\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUHZ0Z2\
        );

    \I__2973\ : InMux
    port map (
            O => \N__13948\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__13945\,
            I => \N__13942\
        );

    \I__2971\ : InMux
    port map (
            O => \N__13942\,
            I => \N__13939\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__13939\,
            I => \N__13936\
        );

    \I__2969\ : Odrv12
    port map (
            O => \N__13936\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIVZ0Z6153\
        );

    \I__2968\ : InMux
    port map (
            O => \N__13933\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__2967\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13927\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__13927\,
            I => \N__13924\
        );

    \I__2965\ : Odrv12
    port map (
            O => \N__13924\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8
        );

    \I__2964\ : InMux
    port map (
            O => \N__13921\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__2963\ : InMux
    port map (
            O => \N__13918\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__13915\,
            I => \N__13912\
        );

    \I__2961\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13905\
        );

    \I__2960\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13905\
        );

    \I__2959\ : InMux
    port map (
            O => \N__13910\,
            I => \N__13902\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__13905\,
            I => \N__13899\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__13902\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3\
        );

    \I__2956\ : Odrv12
    port map (
            O => \N__13899\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3\
        );

    \I__2955\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__13891\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i
        );

    \I__2953\ : InMux
    port map (
            O => \N__13888\,
            I => \N__13882\
        );

    \I__2952\ : InMux
    port map (
            O => \N__13887\,
            I => \N__13877\
        );

    \I__2951\ : InMux
    port map (
            O => \N__13886\,
            I => \N__13877\
        );

    \I__2950\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13873\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__13882\,
            I => \N__13869\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__13877\,
            I => \N__13865\
        );

    \I__2947\ : InMux
    port map (
            O => \N__13876\,
            I => \N__13862\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__13873\,
            I => \N__13859\
        );

    \I__2945\ : InMux
    port map (
            O => \N__13872\,
            I => \N__13855\
        );

    \I__2944\ : Span4Mux_h
    port map (
            O => \N__13869\,
            I => \N__13852\
        );

    \I__2943\ : InMux
    port map (
            O => \N__13868\,
            I => \N__13849\
        );

    \I__2942\ : Span4Mux_h
    port map (
            O => \N__13865\,
            I => \N__13842\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__13862\,
            I => \N__13842\
        );

    \I__2940\ : Span4Mux_h
    port map (
            O => \N__13859\,
            I => \N__13842\
        );

    \I__2939\ : InMux
    port map (
            O => \N__13858\,
            I => \N__13839\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__13855\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__13852\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__13849\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__13842\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__13839\,
            I => charx_if_generate_plus_mult1_un40_sum
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__13828\,
            I => \N__13825\
        );

    \I__2932\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13822\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__13822\,
            I => un5_visiblex_i_0_25
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__13819\,
            I => \N__13816\
        );

    \I__2929\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13813\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__13813\,
            I => column_1_if_generate_plus_mult1_un47_sum1_2
        );

    \I__2927\ : InMux
    port map (
            O => \N__13810\,
            I => column_1_if_generate_plus_mult1_un47_sum_1_cry_1
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__13807\,
            I => \N__13804\
        );

    \I__2925\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13801\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__13801\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\
        );

    \I__2923\ : InMux
    port map (
            O => \N__13798\,
            I => \N__13795\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__13795\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8TZ0Z77\
        );

    \I__2921\ : InMux
    port map (
            O => \N__13792\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__13789\,
            I => \N__13786\
        );

    \I__2919\ : InMux
    port map (
            O => \N__13786\,
            I => \N__13783\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__13783\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0\
        );

    \I__2917\ : InMux
    port map (
            O => \N__13780\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__13777\,
            I => \N__13773\
        );

    \I__2915\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13770\
        );

    \I__2914\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13767\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__13770\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__13767\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf
        );

    \I__2911\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13759\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__13759\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\
        );

    \I__2909\ : InMux
    port map (
            O => \N__13756\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3
        );

    \I__2908\ : InMux
    port map (
            O => \N__13753\,
            I => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4
        );

    \I__2907\ : InMux
    port map (
            O => \N__13750\,
            I => \N__13741\
        );

    \I__2906\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13741\
        );

    \I__2905\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13741\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__13741\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__13738\,
            I => \N__13735\
        );

    \I__2902\ : InMux
    port map (
            O => \N__13735\,
            I => \N__13732\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__13732\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77Z0Z_0\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__13729\,
            I => \N__13726\
        );

    \I__2899\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13723\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__13723\,
            I => charx_i_23
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__13720\,
            I => \N__13716\
        );

    \I__2896\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13710\
        );

    \I__2895\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13705\
        );

    \I__2894\ : InMux
    port map (
            O => \N__13715\,
            I => \N__13705\
        );

    \I__2893\ : InMux
    port map (
            O => \N__13714\,
            I => \N__13702\
        );

    \I__2892\ : InMux
    port map (
            O => \N__13713\,
            I => \N__13699\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__13710\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__13705\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__13702\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__13699\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__13690\,
            I => \N__13685\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__13689\,
            I => \N__13682\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__13688\,
            I => \N__13679\
        );

    \I__2884\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13676\
        );

    \I__2883\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13673\
        );

    \I__2882\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13670\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__13676\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__13673\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__13670\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2\
        );

    \I__2878\ : InMux
    port map (
            O => \N__13663\,
            I => \N__13660\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__13660\,
            I => \N__13653\
        );

    \I__2876\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13650\
        );

    \I__2875\ : InMux
    port map (
            O => \N__13658\,
            I => \N__13645\
        );

    \I__2874\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13645\
        );

    \I__2873\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13642\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__13653\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__13650\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__13645\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__13642\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__13633\,
            I => \N__13630\
        );

    \I__2867\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13627\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__13627\,
            I => charx_i_24
        );

    \I__2865\ : InMux
    port map (
            O => \N__13624\,
            I => \N__13621\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__13621\,
            I => un116_pixel_2_bm_0
        );

    \I__2863\ : InMux
    port map (
            O => \N__13618\,
            I => \N__13615\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__13615\,
            I => \un114_pixel_1_0_3__un116_pixel_5_ns_1_0Z0Z_0\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__13612\,
            I => \N__13608\
        );

    \I__2860\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13604\
        );

    \I__2859\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13600\
        );

    \I__2858\ : InMux
    port map (
            O => \N__13607\,
            I => \N__13596\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__13604\,
            I => \N__13593\
        );

    \I__2856\ : InMux
    port map (
            O => \N__13603\,
            I => \N__13590\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__13600\,
            I => \N__13587\
        );

    \I__2854\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13584\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__13596\,
            I => \N__13581\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__13593\,
            I => \N__13578\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13575\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__13587\,
            I => \N__13572\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__13584\,
            I => \N__13569\
        );

    \I__2848\ : Span4Mux_v
    port map (
            O => \N__13581\,
            I => \N__13564\
        );

    \I__2847\ : Span4Mux_s3_h
    port map (
            O => \N__13578\,
            I => \N__13564\
        );

    \I__2846\ : Span4Mux_s3_v
    port map (
            O => \N__13575\,
            I => \N__13561\
        );

    \I__2845\ : Odrv4
    port map (
            O => \N__13572\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__13569\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__13564\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__13561\,
            I => chessboardpixel_un152_pixel_24
        );

    \I__2841\ : InMux
    port map (
            O => \N__13552\,
            I => \N__13549\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__13549\,
            I => \N__13546\
        );

    \I__2839\ : Odrv4
    port map (
            O => \N__13546\,
            I => \un114_pixel_1_0_3__un116_pixel_6_1_1Z0Z_1\
        );

    \I__2838\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13537\
        );

    \I__2837\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13533\
        );

    \I__2836\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13528\
        );

    \I__2835\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13528\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__13537\,
            I => \N__13525\
        );

    \I__2833\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13522\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__13533\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__13528\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__13525\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__13522\,
            I => charx_if_generate_plus_mult1_un1_sum_axb1
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__13513\,
            I => \N__13510\
        );

    \I__2827\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13506\
        );

    \I__2826\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13503\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__13506\,
            I => \N__13500\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__13503\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4\
        );

    \I__2823\ : Odrv4
    port map (
            O => \N__13500\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4\
        );

    \I__2822\ : InMux
    port map (
            O => \N__13495\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1
        );

    \I__2821\ : InMux
    port map (
            O => \N__13492\,
            I => \N__13489\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__13489\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3EZ0Z987\
        );

    \I__2819\ : InMux
    port map (
            O => \N__13486\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__13483\,
            I => \N__13479\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__13482\,
            I => \N__13476\
        );

    \I__2816\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13471\
        );

    \I__2815\ : InMux
    port map (
            O => \N__13476\,
            I => \N__13471\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__13471\,
            I => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\
        );

    \I__2813\ : InMux
    port map (
            O => \N__13468\,
            I => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__13465\,
            I => \N__13461\
        );

    \I__2811\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13455\
        );

    \I__2810\ : InMux
    port map (
            O => \N__13461\,
            I => \N__13452\
        );

    \I__2809\ : InMux
    port map (
            O => \N__13460\,
            I => \N__13449\
        );

    \I__2808\ : InMux
    port map (
            O => \N__13459\,
            I => \N__13444\
        );

    \I__2807\ : InMux
    port map (
            O => \N__13458\,
            I => \N__13444\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__13455\,
            I => \N__13441\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__13452\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__13449\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__13444\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__13441\,
            I => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987\
        );

    \I__2801\ : InMux
    port map (
            O => \N__13432\,
            I => \N__13429\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__13429\,
            I => un116_pixel_4_am_1
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__13426\,
            I => \N__13419\
        );

    \I__2798\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13414\
        );

    \I__2797\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13409\
        );

    \I__2796\ : InMux
    port map (
            O => \N__13423\,
            I => \N__13409\
        );

    \I__2795\ : InMux
    port map (
            O => \N__13422\,
            I => \N__13406\
        );

    \I__2794\ : InMux
    port map (
            O => \N__13419\,
            I => \N__13403\
        );

    \I__2793\ : InMux
    port map (
            O => \N__13418\,
            I => \N__13400\
        );

    \I__2792\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13397\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__13414\,
            I => \N__13394\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__13409\,
            I => \N_36\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__13406\,
            I => \N_36\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__13403\,
            I => \N_36\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__13400\,
            I => \N_36\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__13397\,
            I => \N_36\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__13394\,
            I => \N_36\
        );

    \I__2784\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13378\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__13378\,
            I => \un116_pixel_5_amZ0Z_5\
        );

    \I__2782\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13372\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__13372\,
            I => \un116_pixel_2_amZ0Z_5\
        );

    \I__2780\ : InMux
    port map (
            O => \N__13369\,
            I => \N__13366\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__13366\,
            I => \N_385\
        );

    \I__2778\ : InMux
    port map (
            O => \N__13363\,
            I => \N__13359\
        );

    \I__2777\ : InMux
    port map (
            O => \N__13362\,
            I => \N__13356\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__13359\,
            I => \N_325\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__13356\,
            I => \N_325\
        );

    \I__2774\ : InMux
    port map (
            O => \N__13351\,
            I => \N__13348\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__13348\,
            I => \un116_pixel_2_bmZ0Z_1\
        );

    \I__2772\ : InMux
    port map (
            O => \N__13345\,
            I => \N__13342\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__13342\,
            I => \un114_pixel_1_0_3__un116_pixel_6_1Z0Z_1\
        );

    \I__2770\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13336\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__13336\,
            I => \N__13331\
        );

    \I__2768\ : InMux
    port map (
            O => \N__13335\,
            I => \N__13328\
        );

    \I__2767\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13325\
        );

    \I__2766\ : Odrv4
    port map (
            O => \N__13331\,
            I => un116_pixel_1_4
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__13328\,
            I => un116_pixel_1_4
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__13325\,
            I => un116_pixel_1_4
        );

    \I__2763\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13314\
        );

    \I__2762\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13311\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__13314\,
            I => \N_374_0\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__13311\,
            I => \N_374_0\
        );

    \I__2759\ : CascadeMux
    port map (
            O => \N__13306\,
            I => \N__13296\
        );

    \I__2758\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13285\
        );

    \I__2757\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13285\
        );

    \I__2756\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13285\
        );

    \I__2755\ : InMux
    port map (
            O => \N__13302\,
            I => \N__13282\
        );

    \I__2754\ : InMux
    port map (
            O => \N__13301\,
            I => \N__13275\
        );

    \I__2753\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13275\
        );

    \I__2752\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13275\
        );

    \I__2751\ : InMux
    port map (
            O => \N__13296\,
            I => \N__13270\
        );

    \I__2750\ : InMux
    port map (
            O => \N__13295\,
            I => \N__13270\
        );

    \I__2749\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13267\
        );

    \I__2748\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13262\
        );

    \I__2747\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13262\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__13285\,
            I => font_un3_pixel_29
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__13282\,
            I => font_un3_pixel_29
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__13275\,
            I => font_un3_pixel_29
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__13270\,
            I => font_un3_pixel_29
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__13267\,
            I => font_un3_pixel_29
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__13262\,
            I => font_un3_pixel_29
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__13249\,
            I => \un116_pixel_7_x0_0_cascade_\
        );

    \I__2739\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13243\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__13243\,
            I => un116_pixel_7_x1_0
        );

    \I__2737\ : InMux
    port map (
            O => \N__13240\,
            I => \N__13237\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__13237\,
            I => un116_pixel_7_ns_0
        );

    \I__2735\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__13231\,
            I => column_0111_0
        );

    \I__2733\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__13225\,
            I => un116_pixel_3_ns_1_0_3
        );

    \I__2731\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13219\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__13219\,
            I => \un114_pixel_1_0_3__g1Z0Z_4\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__13216\,
            I => \N_1583_0_cascade_\
        );

    \I__2728\ : InMux
    port map (
            O => \N__13213\,
            I => \N__13210\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__13210\,
            I => \N_26_0_0\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__13207\,
            I => \un116_pixel_2_amZ0Z_1_cascade_\
        );

    \I__2725\ : InMux
    port map (
            O => \N__13204\,
            I => \N__13201\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__13201\,
            I => un116_pixel_6_1
        );

    \I__2723\ : CascadeMux
    port map (
            O => \N__13198\,
            I => \column_0001_0_cascade_\
        );

    \I__2722\ : InMux
    port map (
            O => \N__13195\,
            I => \N__13192\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__13192\,
            I => \beamY_RNILBST4T2Z0Z_1\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__13189\,
            I => \beamY_RNIT81CMJ2Z0Z_1_cascade_\
        );

    \I__2719\ : InMux
    port map (
            O => \N__13186\,
            I => \N__13183\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__13183\,
            I => \N__13180\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__13180\,
            I => font_un126_pixel_2_am
        );

    \I__2716\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13174\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__13174\,
            I => \N__13171\
        );

    \I__2714\ : Span4Mux_h
    port map (
            O => \N__13171\,
            I => \N__13168\
        );

    \I__2713\ : Odrv4
    port map (
            O => \N__13168\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5RZ0\
        );

    \I__2712\ : InMux
    port map (
            O => \N__13165\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__2711\ : InMux
    port map (
            O => \N__13162\,
            I => \N__13158\
        );

    \I__2710\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13155\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__13158\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__13155\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__13150\,
            I => \N__13147\
        );

    \I__2706\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13144\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__13144\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRDZ0\
        );

    \I__2704\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13138\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__13138\,
            I => \N__13135\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__13135\,
            I => \N__13132\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__13132\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BVZ0Z81\
        );

    \I__2700\ : InMux
    port map (
            O => \N__13129\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__2699\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13123\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__13123\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0LZ0\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__13120\,
            I => \N__13116\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__13119\,
            I => \N__13113\
        );

    \I__2695\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13108\
        );

    \I__2694\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13108\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__13108\,
            I => charx_if_generate_plus_mult1_un61_sum_i_5
        );

    \I__2692\ : InMux
    port map (
            O => \N__13105\,
            I => \N__13102\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__13102\,
            I => \N__13099\
        );

    \I__2690\ : Span4Mux_h
    port map (
            O => \N__13099\,
            I => \N__13096\
        );

    \I__2689\ : Odrv4
    port map (
            O => \N__13096\,
            I => charx_if_generate_plus_mult1_un75_sum_axb_5
        );

    \I__2688\ : InMux
    port map (
            O => \N__13093\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__2687\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13087\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__13087\,
            I => charx_if_generate_plus_mult1_un68_sum_axb_5
        );

    \I__2685\ : InMux
    port map (
            O => \N__13084\,
            I => charx_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__13081\,
            I => \N__13078\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13078\,
            I => \N__13071\
        );

    \I__2682\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13071\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13067\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__13071\,
            I => \N__13064\
        );

    \I__2679\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13061\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__13067\,
            I => \N__13056\
        );

    \I__2677\ : Span4Mux_h
    port map (
            O => \N__13064\,
            I => \N__13056\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__13061\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1\
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__13056\,
            I => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13051\,
            I => \N__13048\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__13048\,
            I => charx_if_generate_plus_mult1_un61_sum_i
        );

    \I__2672\ : InMux
    port map (
            O => \N__13045\,
            I => \N__13042\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__13042\,
            I => \N_41_0\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__13039\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axb_2_sxZ0_cascade_\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__13036\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2_cascade_\
        );

    \I__2668\ : InMux
    port map (
            O => \N__13033\,
            I => \N__13030\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__13030\,
            I => if_generate_plus_mult1_un54_sum_axb_2_l_fx
        );

    \I__2666\ : InMux
    port map (
            O => \N__13027\,
            I => \N__13024\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__13024\,
            I => column_1_if_generate_plus_mult1_un47_sum0_4
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__13021\,
            I => \if_generate_plus_mult1_un47_sum_m_5_cascade_\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13018\,
            I => \N__13015\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__13015\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\
        );

    \I__2661\ : InMux
    port map (
            O => \N__13012\,
            I => \N__13009\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__13009\,
            I => column_1_if_generate_plus_mult1_un47_sum0_2
        );

    \I__2659\ : InMux
    port map (
            O => \N__13006\,
            I => \N__13001\
        );

    \I__2658\ : InMux
    port map (
            O => \N__13005\,
            I => \N__12996\
        );

    \I__2657\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12996\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__13001\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__12996\,
            I => if_generate_plus_mult1_un47_sum_m_5
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__12991\,
            I => \N__12988\
        );

    \I__2653\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12985\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__12985\,
            I => if_generate_plus_mult1_un54_sum_axb_3_l_fx
        );

    \I__2651\ : InMux
    port map (
            O => \N__12982\,
            I => \N__12976\
        );

    \I__2650\ : InMux
    port map (
            O => \N__12981\,
            I => \N__12969\
        );

    \I__2649\ : InMux
    port map (
            O => \N__12980\,
            I => \N__12969\
        );

    \I__2648\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12969\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__12976\,
            I => column_1_if_generate_plus_mult1_un47_sum0_5
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__12969\,
            I => column_1_if_generate_plus_mult1_un47_sum0_5
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__12964\,
            I => \N__12960\
        );

    \I__2644\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \N__12957\
        );

    \I__2643\ : InMux
    port map (
            O => \N__12960\,
            I => \N__12950\
        );

    \I__2642\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12950\
        );

    \I__2641\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12947\
        );

    \I__2640\ : InMux
    port map (
            O => \N__12955\,
            I => \N__12944\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__12950\,
            I => \N_584_i\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__12947\,
            I => \N_584_i\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__12944\,
            I => \N_584_i\
        );

    \I__2636\ : InMux
    port map (
            O => \N__12937\,
            I => \N__12931\
        );

    \I__2635\ : InMux
    port map (
            O => \N__12936\,
            I => \N__12928\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__12935\,
            I => \N__12925\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__12934\,
            I => \N__12920\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__12931\,
            I => \N__12915\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__12928\,
            I => \N__12912\
        );

    \I__2630\ : InMux
    port map (
            O => \N__12925\,
            I => \N__12907\
        );

    \I__2629\ : InMux
    port map (
            O => \N__12924\,
            I => \N__12907\
        );

    \I__2628\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12902\
        );

    \I__2627\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12902\
        );

    \I__2626\ : InMux
    port map (
            O => \N__12919\,
            I => \N__12897\
        );

    \I__2625\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12897\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__12915\,
            I => \N__12885\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__12912\,
            I => \N__12885\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__12907\,
            I => \N__12885\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__12902\,
            I => \N__12885\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__12897\,
            I => \N__12885\
        );

    \I__2619\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12882\
        );

    \I__2618\ : Odrv4
    port map (
            O => \N__12885\,
            I => \N_37_i\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__12882\,
            I => \N_37_i\
        );

    \I__2616\ : InMux
    port map (
            O => \N__12877\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__12874\,
            I => \N__12871\
        );

    \I__2614\ : InMux
    port map (
            O => \N__12871\,
            I => \N__12868\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__12868\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_invZ0\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12865\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__12862\,
            I => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843_cascade_\
        );

    \I__2610\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12856\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__12856\,
            I => charx_if_generate_plus_mult1_un68_sum_i
        );

    \I__2608\ : CascadeMux
    port map (
            O => \N__12853\,
            I => \N__12850\
        );

    \I__2607\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12847\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__12847\,
            I => \N__12844\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__12844\,
            I => \un114_pixel_1_0_3__un4_row_8Z0Z_0\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__12841\,
            I => \N__12838\
        );

    \I__2603\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12835\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__12835\,
            I => charx_if_generate_plus_mult1_un68_sum_i_5
        );

    \I__2601\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12829\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__12829\,
            I => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx
        );

    \I__2599\ : InMux
    port map (
            O => \N__12826\,
            I => \N__12823\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__12823\,
            I => \un114_pixel_1_0_3__font_un57_pixelZ0Z_0\
        );

    \I__2597\ : InMux
    port map (
            O => \N__12820\,
            I => \N__12817\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__12817\,
            I => \N__12813\
        );

    \I__2595\ : InMux
    port map (
            O => \N__12816\,
            I => \N__12806\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__12813\,
            I => \N__12801\
        );

    \I__2593\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12798\
        );

    \I__2592\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12793\
        );

    \I__2591\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12793\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__12809\,
            I => \N__12788\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__12806\,
            I => \N__12785\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12782\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__12804\,
            I => \N__12779\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__12801\,
            I => \N__12772\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__12798\,
            I => \N__12772\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__12793\,
            I => \N__12772\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12769\
        );

    \I__2582\ : InMux
    port map (
            O => \N__12791\,
            I => \N__12766\
        );

    \I__2581\ : InMux
    port map (
            O => \N__12788\,
            I => \N__12763\
        );

    \I__2580\ : Span4Mux_h
    port map (
            O => \N__12785\,
            I => \N__12758\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__12782\,
            I => \N__12758\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12755\
        );

    \I__2577\ : Span4Mux_v
    port map (
            O => \N__12772\,
            I => \N__12752\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__12769\,
            I => \N__12749\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__12766\,
            I => \N__12744\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__12763\,
            I => \N__12744\
        );

    \I__2573\ : Span4Mux_v
    port map (
            O => \N__12758\,
            I => \N__12739\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__12755\,
            I => \N__12739\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__12752\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__12749\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2569\ : Odrv12
    port map (
            O => \N__12744\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2568\ : Odrv4
    port map (
            O => \N__12739\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum
        );

    \I__2567\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12727\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__12727\,
            I => \N__12724\
        );

    \I__2565\ : Span4Mux_h
    port map (
            O => \N__12724\,
            I => \N__12718\
        );

    \I__2564\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12715\
        );

    \I__2563\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12710\
        );

    \I__2562\ : InMux
    port map (
            O => \N__12721\,
            I => \N__12710\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__12718\,
            I => if_generate_plus_mult1_un61_sum_axbxc5
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__12715\,
            I => if_generate_plus_mult1_un61_sum_axbxc5
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__12710\,
            I => if_generate_plus_mult1_un61_sum_axbxc5
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__12703\,
            I => \un114_pixel_1_0_3__un4_row_8Z0Z_3_cascade_\
        );

    \I__2557\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12697\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__12697\,
            I => \N__12694\
        );

    \I__2555\ : Odrv4
    port map (
            O => \N__12694\,
            I => \un114_pixel_1_0_3__un4_row_8_7Z0Z_1\
        );

    \I__2554\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12680\
        );

    \I__2553\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12680\
        );

    \I__2552\ : InMux
    port map (
            O => \N__12689\,
            I => \N__12674\
        );

    \I__2551\ : InMux
    port map (
            O => \N__12688\,
            I => \N__12674\
        );

    \I__2550\ : InMux
    port map (
            O => \N__12687\,
            I => \N__12671\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__12686\,
            I => \N__12667\
        );

    \I__2548\ : CascadeMux
    port map (
            O => \N__12685\,
            I => \N__12662\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__12680\,
            I => \N__12659\
        );

    \I__2546\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12656\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__12674\,
            I => \N__12651\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__12671\,
            I => \N__12648\
        );

    \I__2543\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12641\
        );

    \I__2542\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12641\
        );

    \I__2541\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12641\
        );

    \I__2540\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12636\
        );

    \I__2539\ : InMux
    port map (
            O => \N__12662\,
            I => \N__12636\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__12659\,
            I => \N__12631\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__12656\,
            I => \N__12631\
        );

    \I__2536\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12626\
        );

    \I__2535\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12626\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__12651\,
            I => \N__12623\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__12648\,
            I => \N__12620\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__12641\,
            I => \N__12615\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__12636\,
            I => \N__12615\
        );

    \I__2530\ : Span4Mux_h
    port map (
            O => \N__12631\,
            I => \N__12610\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__12626\,
            I => \N__12610\
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__12623\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum
        );

    \I__2527\ : Odrv4
    port map (
            O => \N__12620\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__12615\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum
        );

    \I__2525\ : Odrv4
    port map (
            O => \N__12610\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum
        );

    \I__2524\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12593\
        );

    \I__2523\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12593\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__12599\,
            I => \N__12588\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__12598\,
            I => \N__12585\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__12593\,
            I => \N__12578\
        );

    \I__2519\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12575\
        );

    \I__2518\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12572\
        );

    \I__2517\ : InMux
    port map (
            O => \N__12588\,
            I => \N__12567\
        );

    \I__2516\ : InMux
    port map (
            O => \N__12585\,
            I => \N__12567\
        );

    \I__2515\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12560\
        );

    \I__2514\ : InMux
    port map (
            O => \N__12583\,
            I => \N__12560\
        );

    \I__2513\ : InMux
    port map (
            O => \N__12582\,
            I => \N__12560\
        );

    \I__2512\ : InMux
    port map (
            O => \N__12581\,
            I => \N__12557\
        );

    \I__2511\ : Span4Mux_v
    port map (
            O => \N__12578\,
            I => \N__12554\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__12575\,
            I => \N__12551\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__12572\,
            I => \N__12548\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__12567\,
            I => \N__12545\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__12560\,
            I => \N__12540\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__12557\,
            I => \N__12540\
        );

    \I__2505\ : Span4Mux_h
    port map (
            O => \N__12554\,
            I => \N__12533\
        );

    \I__2504\ : Span4Mux_v
    port map (
            O => \N__12551\,
            I => \N__12533\
        );

    \I__2503\ : Span4Mux_h
    port map (
            O => \N__12548\,
            I => \N__12530\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__12545\,
            I => \N__12525\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__12540\,
            I => \N__12525\
        );

    \I__2500\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12522\
        );

    \I__2499\ : InMux
    port map (
            O => \N__12538\,
            I => \N__12519\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__12533\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__12530\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__12525\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__12522\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__12519\,
            I => chary_if_generate_plus_mult1_un33_sum_axb3
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__12508\,
            I => \N__12504\
        );

    \I__2492\ : InMux
    port map (
            O => \N__12507\,
            I => \N__12500\
        );

    \I__2491\ : InMux
    port map (
            O => \N__12504\,
            I => \N__12494\
        );

    \I__2490\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12494\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12500\,
            I => \N__12491\
        );

    \I__2488\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12488\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__12494\,
            I => \N__12485\
        );

    \I__2486\ : Odrv4
    port map (
            O => \N__12491\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__12488\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__2484\ : Odrv12
    port map (
            O => \N__12485\,
            I => if_generate_plus_mult1_un54_sum_s_5
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__12478\,
            I => \N__12475\
        );

    \I__2482\ : InMux
    port map (
            O => \N__12475\,
            I => \N__12472\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__12472\,
            I => \un114_pixel_1_0_3__un4_row_8Z0Z_2\
        );

    \I__2480\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12466\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__12466\,
            I => \N__12462\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__12465\,
            I => \N__12459\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__12462\,
            I => \N__12456\
        );

    \I__2476\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12453\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__12456\,
            I => \row_1_if_generate_plus_mult1_un75_sum_cZ0Z5\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__12453\,
            I => \row_1_if_generate_plus_mult1_un75_sum_cZ0Z5\
        );

    \I__2473\ : InMux
    port map (
            O => \N__12448\,
            I => \N__12442\
        );

    \I__2472\ : InMux
    port map (
            O => \N__12447\,
            I => \N__12442\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12439\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__12439\,
            I => \N__12433\
        );

    \I__2469\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12430\
        );

    \I__2468\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12425\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12436\,
            I => \N__12425\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__12433\,
            I => if_generate_plus_mult1_un68_sum_axbxc5
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__12430\,
            I => if_generate_plus_mult1_un68_sum_axbxc5
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__12425\,
            I => if_generate_plus_mult1_un68_sum_axbxc5
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__12418\,
            I => \N__12414\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__12417\,
            I => \N__12411\
        );

    \I__2461\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12407\
        );

    \I__2460\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12401\
        );

    \I__2459\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12401\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12398\
        );

    \I__2457\ : InMux
    port map (
            O => \N__12406\,
            I => \N__12395\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__12401\,
            I => \N__12392\
        );

    \I__2455\ : Span4Mux_h
    port map (
            O => \N__12398\,
            I => \N__12389\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__12395\,
            I => \N__12386\
        );

    \I__2453\ : Span4Mux_h
    port map (
            O => \N__12392\,
            I => \N__12383\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__12389\,
            I => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__12386\,
            I => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__12383\,
            I => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2\
        );

    \I__2449\ : InMux
    port map (
            O => \N__12376\,
            I => \N__12373\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__12373\,
            I => \un114_pixel_1_0_3__un4_row_8Z0Z_7\
        );

    \I__2447\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12367\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__12367\,
            I => \un114_pixel_1_0_3__un4_rowZ0Z_8\
        );

    \I__2445\ : InMux
    port map (
            O => \N__12364\,
            I => \N__12361\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__12361\,
            I => \N__12357\
        );

    \I__2443\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12354\
        );

    \I__2442\ : Span4Mux_h
    port map (
            O => \N__12357\,
            I => \N__12351\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__12354\,
            I => \N__12348\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__12351\,
            I => \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1\
        );

    \I__2439\ : Odrv12
    port map (
            O => \N__12348\,
            I => \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1\
        );

    \I__2438\ : InMux
    port map (
            O => \N__12343\,
            I => \N__12339\
        );

    \I__2437\ : InMux
    port map (
            O => \N__12342\,
            I => \N__12336\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__12339\,
            I => \N__12333\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__12336\,
            I => \N__12330\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__12333\,
            I => \N__12325\
        );

    \I__2433\ : Span4Mux_h
    port map (
            O => \N__12330\,
            I => \N__12325\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__12325\,
            I => row_1_if_generate_plus_mult1_un82_sum_c5
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__12322\,
            I => \un114_pixel_1_0_3__un4_rowZ0Z_8_cascade_\
        );

    \I__2430\ : InMux
    port map (
            O => \N__12319\,
            I => \N__12316\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__12316\,
            I => \N__12313\
        );

    \I__2428\ : Odrv12
    port map (
            O => \N__12313\,
            I => \un114_pixel_1_0_3__Pixel_3_sqmuxaZ0Z_0\
        );

    \I__2427\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12307\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__12307\,
            I => \N__12303\
        );

    \I__2425\ : InMux
    port map (
            O => \N__12306\,
            I => \N__12300\
        );

    \I__2424\ : Odrv4
    port map (
            O => \N__12303\,
            I => \Pixel_3_sqmuxa\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__12300\,
            I => \Pixel_3_sqmuxa\
        );

    \I__2422\ : InMux
    port map (
            O => \N__12295\,
            I => charx_if_generate_plus_mult1_un75_sum_cry_1
        );

    \I__2421\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12288\
        );

    \I__2420\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12285\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__12288\,
            I => \N__12282\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__12285\,
            I => \N__12275\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__12282\,
            I => \N__12275\
        );

    \I__2416\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12270\
        );

    \I__2415\ : InMux
    port map (
            O => \N__12280\,
            I => \N__12270\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__12275\,
            I => \beamY_RNIHHB5F01Z0Z_4\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__12270\,
            I => \beamY_RNIHHB5F01Z0Z_4\
        );

    \I__2412\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12260\
        );

    \I__2411\ : InMux
    port map (
            O => \N__12264\,
            I => \N__12255\
        );

    \I__2410\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12255\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__12260\,
            I => \N__12242\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__12255\,
            I => \N__12239\
        );

    \I__2407\ : InMux
    port map (
            O => \N__12254\,
            I => \N__12234\
        );

    \I__2406\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12234\
        );

    \I__2405\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12231\
        );

    \I__2404\ : InMux
    port map (
            O => \N__12251\,
            I => \N__12228\
        );

    \I__2403\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12225\
        );

    \I__2402\ : InMux
    port map (
            O => \N__12249\,
            I => \N__12222\
        );

    \I__2401\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12217\
        );

    \I__2400\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12217\
        );

    \I__2399\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12212\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12209\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__12242\,
            I => \N__12203\
        );

    \I__2396\ : Span4Mux_v
    port map (
            O => \N__12239\,
            I => \N__12203\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__12234\,
            I => \N__12196\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__12231\,
            I => \N__12196\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__12228\,
            I => \N__12196\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__12225\,
            I => \N__12189\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__12222\,
            I => \N__12189\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__12217\,
            I => \N__12189\
        );

    \I__2389\ : InMux
    port map (
            O => \N__12216\,
            I => \N__12184\
        );

    \I__2388\ : InMux
    port map (
            O => \N__12215\,
            I => \N__12184\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__12212\,
            I => \N__12179\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__12209\,
            I => \N__12179\
        );

    \I__2385\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12174\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__12203\,
            I => \N__12171\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__12196\,
            I => \N__12164\
        );

    \I__2382\ : Span4Mux_v
    port map (
            O => \N__12189\,
            I => \N__12164\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__12184\,
            I => \N__12164\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__12179\,
            I => \N__12161\
        );

    \I__2379\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12156\
        );

    \I__2378\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12156\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__12174\,
            I => \beamYZ0Z_2\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__12171\,
            I => \beamYZ0Z_2\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__12164\,
            I => \beamYZ0Z_2\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__12161\,
            I => \beamYZ0Z_2\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__12156\,
            I => \beamYZ0Z_2\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__12145\,
            I => \N__12142\
        );

    \I__2371\ : InMux
    port map (
            O => \N__12142\,
            I => \N__12139\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__12139\,
            I => \beamY_RNI7OE17CZ0Z_0\
        );

    \I__2369\ : InMux
    port map (
            O => \N__12136\,
            I => \N__12133\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__12133\,
            I => \N__12130\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__12130\,
            I => \beamY_RNIVU1O9RZ0Z_1\
        );

    \I__2366\ : InMux
    port map (
            O => \N__12127\,
            I => \N__12124\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__12124\,
            I => font_un126_pixel_6_bm
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__12121\,
            I => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\
        );

    \I__2363\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12114\
        );

    \I__2362\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12111\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__12114\,
            I => \N__12108\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__12111\,
            I => \N__12105\
        );

    \I__2359\ : Span4Mux_v
    port map (
            O => \N__12108\,
            I => \N__12102\
        );

    \I__2358\ : Span4Mux_h
    port map (
            O => \N__12105\,
            I => \N__12099\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__12102\,
            I => un15_beamy
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__12099\,
            I => un15_beamy
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__12094\,
            I => \r_i1_mux_cascade_\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__12091\,
            I => \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_1_cascade_\
        );

    \I__2353\ : InMux
    port map (
            O => \N__12088\,
            I => \N__12085\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__12085\,
            I => \N__12082\
        );

    \I__2351\ : Span4Mux_v
    port map (
            O => \N__12082\,
            I => \N__12079\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__12079\,
            I => chary_24
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__12076\,
            I => \un114_pixel_1_0_3__font_un126_pixel_m_1_0_cascade_\
        );

    \I__2348\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12070\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__12070\,
            I => chary_23
        );

    \I__2346\ : InMux
    port map (
            O => \N__12067\,
            I => \N__12064\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__12064\,
            I => \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3\
        );

    \I__2344\ : InMux
    port map (
            O => \N__12061\,
            I => \N__12057\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12054\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__12057\,
            I => \N__12051\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__12054\,
            I => \N__12048\
        );

    \I__2340\ : Span4Mux_h
    port map (
            O => \N__12051\,
            I => \N__12045\
        );

    \I__2339\ : Span12Mux_s5_v
    port map (
            O => \N__12048\,
            I => \N__12042\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__12045\,
            I => \N__12039\
        );

    \I__2337\ : Odrv12
    port map (
            O => \N__12042\,
            I => un1_beamylto9
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__12039\,
            I => un1_beamylto9
        );

    \I__2335\ : CascadeMux
    port map (
            O => \N__12034\,
            I => \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3_cascade_\
        );

    \I__2334\ : InMux
    port map (
            O => \N__12031\,
            I => \N__12028\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__12028\,
            I => \Pixel_r_sn\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__12025\,
            I => \N__12020\
        );

    \I__2331\ : CascadeMux
    port map (
            O => \N__12024\,
            I => \N__12015\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12023\,
            I => \N__12012\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12020\,
            I => \N__12009\
        );

    \I__2328\ : InMux
    port map (
            O => \N__12019\,
            I => \N__12004\
        );

    \I__2327\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12004\
        );

    \I__2326\ : InMux
    port map (
            O => \N__12015\,
            I => \N__11999\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__12012\,
            I => \N__11994\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__12009\,
            I => \N__11994\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12004\,
            I => \N__11991\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__12003\,
            I => \N__11985\
        );

    \I__2321\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11982\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__11999\,
            I => \N__11979\
        );

    \I__2319\ : Span4Mux_h
    port map (
            O => \N__11994\,
            I => \N__11976\
        );

    \I__2318\ : Span4Mux_h
    port map (
            O => \N__11991\,
            I => \N__11973\
        );

    \I__2317\ : InMux
    port map (
            O => \N__11990\,
            I => \N__11966\
        );

    \I__2316\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11966\
        );

    \I__2315\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11966\
        );

    \I__2314\ : InMux
    port map (
            O => \N__11985\,
            I => \N__11963\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__11982\,
            I => \beamXZ0Z_0\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__11979\,
            I => \beamXZ0Z_0\
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__11976\,
            I => \beamXZ0Z_0\
        );

    \I__2310\ : Odrv4
    port map (
            O => \N__11973\,
            I => \beamXZ0Z_0\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__11966\,
            I => \beamXZ0Z_0\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__11963\,
            I => \beamXZ0Z_0\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__11950\,
            I => \N_364_cascade_\
        );

    \I__2306\ : CascadeMux
    port map (
            O => \N__11947\,
            I => \un116_pixel_7_ns_1_4_cascade_\
        );

    \I__2305\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11941\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__11941\,
            I => \beamY_RNI2L0T663Z0Z_0\
        );

    \I__2303\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11935\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__11935\,
            I => column_0111_1_0
        );

    \I__2301\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11929\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__11929\,
            I => \beamY_RNI1J75181Z0Z_1\
        );

    \I__2299\ : CascadeMux
    port map (
            O => \N__11926\,
            I => \font_un126_pixel_6_am_cascade_\
        );

    \I__2298\ : InMux
    port map (
            O => \N__11923\,
            I => \N__11920\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__11920\,
            I => \N__11917\
        );

    \I__2296\ : Span4Mux_h
    port map (
            O => \N__11917\,
            I => \N__11914\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__11914\,
            I => un1_beamy_0
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__11911\,
            I => \N_1075_0_cascade_\
        );

    \I__2293\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11905\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__11905\,
            I => \N__11902\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__11902\,
            I => \N_400\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__11899\,
            I => \Pixel_r_rn_0_cascade_\
        );

    \I__2289\ : IoInMux
    port map (
            O => \N__11896\,
            I => \N__11893\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__11893\,
            I => \N__11890\
        );

    \I__2287\ : Span4Mux_s3_v
    port map (
            O => \N__11890\,
            I => \N__11887\
        );

    \I__2286\ : Odrv4
    port map (
            O => \N__11887\,
            I => \Pixel_c\
        );

    \I__2285\ : ClkMux
    port map (
            O => \N__11884\,
            I => \N__11845\
        );

    \I__2284\ : ClkMux
    port map (
            O => \N__11883\,
            I => \N__11845\
        );

    \I__2283\ : ClkMux
    port map (
            O => \N__11882\,
            I => \N__11845\
        );

    \I__2282\ : ClkMux
    port map (
            O => \N__11881\,
            I => \N__11845\
        );

    \I__2281\ : ClkMux
    port map (
            O => \N__11880\,
            I => \N__11845\
        );

    \I__2280\ : ClkMux
    port map (
            O => \N__11879\,
            I => \N__11845\
        );

    \I__2279\ : ClkMux
    port map (
            O => \N__11878\,
            I => \N__11845\
        );

    \I__2278\ : ClkMux
    port map (
            O => \N__11877\,
            I => \N__11845\
        );

    \I__2277\ : ClkMux
    port map (
            O => \N__11876\,
            I => \N__11845\
        );

    \I__2276\ : ClkMux
    port map (
            O => \N__11875\,
            I => \N__11845\
        );

    \I__2275\ : ClkMux
    port map (
            O => \N__11874\,
            I => \N__11845\
        );

    \I__2274\ : ClkMux
    port map (
            O => \N__11873\,
            I => \N__11845\
        );

    \I__2273\ : ClkMux
    port map (
            O => \N__11872\,
            I => \N__11845\
        );

    \I__2272\ : GlobalMux
    port map (
            O => \N__11845\,
            I => \N__11842\
        );

    \I__2271\ : gio2CtrlBuf
    port map (
            O => \N__11842\,
            I => \PixelClock_g\
        );

    \I__2270\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11836\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__11836\,
            I => \N__11833\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__11833\,
            I => \N__11830\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__11830\,
            I => font_un28_pixel_0_0_29
        );

    \I__2266\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11824\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__11824\,
            I => font_un126_pixel_2_bm
        );

    \I__2264\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11818\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__11818\,
            I => \un114_pixel_1_0_3__font_un126_pixel_7_d_ns_1_0_0\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__11815\,
            I => \font_un3_pixel_29_cascade_\
        );

    \I__2261\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11809\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__11809\,
            I => un116_pixel_5_bm_6
        );

    \I__2259\ : InMux
    port map (
            O => \N__11806\,
            I => \N__11803\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__11803\,
            I => un116_pixel_4_bm_1
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__11800\,
            I => \beamY_RNI1C50FS3Z0Z_0_cascade_\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__11797\,
            I => \un116_pixel_3_bm_1_6_cascade_\
        );

    \I__2255\ : InMux
    port map (
            O => \N__11794\,
            I => \N__11788\
        );

    \I__2254\ : InMux
    port map (
            O => \N__11793\,
            I => \N__11788\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__11788\,
            I => \N__11785\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__11785\,
            I => \beamY_RNIOHI2NGZ0Z_0\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__11782\,
            I => \N_1556_0_cascade_\
        );

    \I__2250\ : InMux
    port map (
            O => \N__11779\,
            I => \N__11776\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__11776\,
            I => \N__11773\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__11773\,
            I => \N_347_0\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__11770\,
            I => \N__11767\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11764\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__11764\,
            I => font_un28_pixel_0_29
        );

    \I__2244\ : InMux
    port map (
            O => \N__11761\,
            I => \N__11758\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__11758\,
            I => \N_368_0\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__11755\,
            I => \un114_pixel_1_0_3__font_un126_pixel_1_d_ns_1_0_cascade_\
        );

    \I__2241\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11749\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__11749\,
            I => \N_389_0\
        );

    \I__2239\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11743\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__11743\,
            I => \N_346_0_0_1\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__11740\,
            I => \g0_cascade_\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__11737\,
            I => \N_36_cascade_\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__11734\,
            I => \un116_pixel_3_ns_1_1_cascade_\
        );

    \I__2234\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11728\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__11728\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLMZ0Z67\
        );

    \I__2232\ : InMux
    port map (
            O => \N__11725\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__2231\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11719\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__11719\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSAZ0\
        );

    \I__2229\ : InMux
    port map (
            O => \N__11716\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__2228\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11710\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__11710\,
            I => charx_if_generate_plus_mult1_un61_sum_axb_5
        );

    \I__2226\ : InMux
    port map (
            O => \N__11707\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__11704\,
            I => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0_cascade_\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__11701\,
            I => \N__11697\
        );

    \I__2223\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11693\
        );

    \I__2222\ : InMux
    port map (
            O => \N__11697\,
            I => \N__11688\
        );

    \I__2221\ : InMux
    port map (
            O => \N__11696\,
            I => \N__11688\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__11693\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__11688\,
            I => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__11683\,
            I => \N__11679\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__11682\,
            I => \N__11676\
        );

    \I__2216\ : InMux
    port map (
            O => \N__11679\,
            I => \N__11671\
        );

    \I__2215\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11671\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__11671\,
            I => charx_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__2213\ : IoInMux
    port map (
            O => \N__11668\,
            I => \N__11665\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__11665\,
            I => \VSync_c\
        );

    \I__2211\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__11659\,
            I => un116_pixel_3_am_2
        );

    \I__2209\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11653\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__11653\,
            I => \N__11646\
        );

    \I__2207\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11642\
        );

    \I__2206\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11637\
        );

    \I__2205\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11637\
        );

    \I__2204\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11634\
        );

    \I__2203\ : Span4Mux_v
    port map (
            O => \N__11646\,
            I => \N__11631\
        );

    \I__2202\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11628\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__11642\,
            I => \N__11623\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__11637\,
            I => \N__11623\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__11634\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__11631\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__11628\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__11623\,
            I => charx_if_generate_plus_mult1_un47_sum
        );

    \I__2195\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11611\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__11611\,
            I => charx_if_generate_plus_mult1_un47_sum_i
        );

    \I__2193\ : InMux
    port map (
            O => \N__11608\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__2192\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11601\
        );

    \I__2191\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11598\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__11601\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__11598\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__11593\,
            I => \N__11590\
        );

    \I__2187\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11587\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__11587\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0OZ0Z3\
        );

    \I__2185\ : InMux
    port map (
            O => \N__11584\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__2184\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11578\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__11578\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCDZ0Z16\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__11575\,
            I => \N__11571\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__11574\,
            I => \N__11568\
        );

    \I__2180\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11563\
        );

    \I__2179\ : InMux
    port map (
            O => \N__11568\,
            I => \N__11563\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__11563\,
            I => charx_if_generate_plus_mult1_un47_sum_i_5
        );

    \I__2177\ : InMux
    port map (
            O => \N__11560\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__2176\ : InMux
    port map (
            O => \N__11557\,
            I => \N__11554\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__11554\,
            I => charx_if_generate_plus_mult1_un54_sum_axb_5
        );

    \I__2174\ : InMux
    port map (
            O => \N__11551\,
            I => charx_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2173\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11539\
        );

    \I__2172\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11539\
        );

    \I__2171\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11532\
        );

    \I__2170\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11532\
        );

    \I__2169\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11529\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__11539\,
            I => \N__11526\
        );

    \I__2167\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11523\
        );

    \I__2166\ : InMux
    port map (
            O => \N__11537\,
            I => \N__11520\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__11532\,
            I => \N__11517\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__11529\,
            I => \N__11514\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__11526\,
            I => \N__11511\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__11523\,
            I => \N__11506\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__11520\,
            I => \N__11506\
        );

    \I__2160\ : Span4Mux_s3_v
    port map (
            O => \N__11517\,
            I => \N__11503\
        );

    \I__2159\ : Odrv12
    port map (
            O => \N__11514\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__11511\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__2157\ : Odrv4
    port map (
            O => \N__11506\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__11503\,
            I => charx_if_generate_plus_mult1_un54_sum
        );

    \I__2155\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11491\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__11491\,
            I => charx_if_generate_plus_mult1_un54_sum_i
        );

    \I__2153\ : InMux
    port map (
            O => \N__11488\,
            I => charx_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__2152\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11482\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__11482\,
            I => column_1_if_generate_plus_mult1_un47_sum0_3
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__11479\,
            I => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_\
        );

    \I__2149\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11473\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__11473\,
            I => if_generate_plus_mult1_un54_sum_axb_4_l_fx
        );

    \I__2147\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11467\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__11467\,
            I => \N__11464\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__11464\,
            I => charx_if_generate_plus_mult1_un40_sum_i
        );

    \I__2144\ : InMux
    port map (
            O => \N__11461\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_1
        );

    \I__2143\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11453\
        );

    \I__2142\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11450\
        );

    \I__2141\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11447\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__11453\,
            I => \N__11442\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__11450\,
            I => \N__11442\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__11447\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__11442\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__2135\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11431\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__2133\ : Odrv12
    port map (
            O => \N__11428\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEBZ0Z2\
        );

    \I__2132\ : InMux
    port map (
            O => \N__11425\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__2131\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11419\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11416\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__11416\,
            I => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLITZ0Z2\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__11413\,
            I => \N__11409\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__11412\,
            I => \N__11406\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11401\
        );

    \I__2125\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11401\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__11401\,
            I => charx_if_generate_plus_mult1_un40_sum_i_5
        );

    \I__2123\ : InMux
    port map (
            O => \N__11398\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__2122\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__11392\,
            I => \N__11389\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__11389\,
            I => charx_if_generate_plus_mult1_un47_sum_axb_5
        );

    \I__2119\ : InMux
    port map (
            O => \N__11386\,
            I => charx_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__11383\,
            I => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6_cascade_\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__11380\,
            I => \N__11377\
        );

    \I__2116\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11374\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__11374\,
            I => un5_visiblex_i_25
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__11371\,
            I => \N__11368\
        );

    \I__2113\ : InMux
    port map (
            O => \N__11368\,
            I => \N__11365\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__11365\,
            I => if_generate_plus_mult1_un47_sum_0_cry_3_ma
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__11362\,
            I => \N__11359\
        );

    \I__2110\ : InMux
    port map (
            O => \N__11359\,
            I => \N__11356\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__11356\,
            I => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx
        );

    \I__2108\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11350\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11347\
        );

    \I__2106\ : Span4Mux_h
    port map (
            O => \N__11347\,
            I => \N__11344\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__11344\,
            I => if_generate_plus_mult1_un54_sum_cry_2_s
        );

    \I__2104\ : InMux
    port map (
            O => \N__11341\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_1
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__11338\,
            I => \N__11335\
        );

    \I__2102\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11332\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__11332\,
            I => \N__11329\
        );

    \I__2100\ : Span4Mux_h
    port map (
            O => \N__11329\,
            I => \N__11326\
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__11326\,
            I => if_generate_plus_mult1_un54_sum_cry_3_s
        );

    \I__2098\ : InMux
    port map (
            O => \N__11323\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__2097\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11317\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__11317\,
            I => \N__11314\
        );

    \I__2095\ : Odrv12
    port map (
            O => \N__11314\,
            I => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\
        );

    \I__2094\ : InMux
    port map (
            O => \N__11311\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__2093\ : InMux
    port map (
            O => \N__11308\,
            I => column_1_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__2092\ : InMux
    port map (
            O => \N__11305\,
            I => \N__11302\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__11302\,
            I => charx_if_generate_plus_mult1_un40_sum_axb_5
        );

    \I__2090\ : InMux
    port map (
            O => \N__11299\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__2089\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__11293\,
            I => charx_if_generate_plus_mult1_un33_sum_i
        );

    \I__2087\ : InMux
    port map (
            O => \N__11290\,
            I => \N__11287\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__11287\,
            I => charx_if_generate_plus_mult1_un26_sum_i
        );

    \I__2085\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11281\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__11281\,
            I => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx
        );

    \I__2083\ : InMux
    port map (
            O => \N__11278\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_1
        );

    \I__2082\ : InMux
    port map (
            O => \N__11275\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_2
        );

    \I__2081\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__11269\,
            I => \N__11266\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__11266\,
            I => \N_204_0_i\
        );

    \I__2078\ : InMux
    port map (
            O => \N__11263\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_3
        );

    \I__2077\ : InMux
    port map (
            O => \N__11260\,
            I => column_1_if_generate_plus_mult1_un47_sum_0_cry_4
        );

    \I__2076\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11254\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__11254\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\
        );

    \I__2074\ : InMux
    port map (
            O => \N__11251\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__2073\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11245\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__11245\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HLZ0\
        );

    \I__2071\ : InMux
    port map (
            O => \N__11242\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__2070\ : InMux
    port map (
            O => \N__11239\,
            I => \N__11236\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__11236\,
            I => charx_if_generate_plus_mult1_un33_sum_axb_5
        );

    \I__2068\ : InMux
    port map (
            O => \N__11233\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__11230\,
            I => \N__11226\
        );

    \I__2066\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11222\
        );

    \I__2065\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11217\
        );

    \I__2064\ : InMux
    port map (
            O => \N__11225\,
            I => \N__11217\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__11222\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__11217\,
            I => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\
        );

    \I__2061\ : CascadeMux
    port map (
            O => \N__11212\,
            I => \N__11208\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__11211\,
            I => \N__11205\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11208\,
            I => \N__11200\
        );

    \I__2058\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11200\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__11200\,
            I => charx_if_generate_plus_mult1_un26_sum_i_5
        );

    \I__2056\ : InMux
    port map (
            O => \N__11197\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_1
        );

    \I__2055\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11189\
        );

    \I__2054\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11186\
        );

    \I__2053\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11183\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__11189\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__11186\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__11183\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__11176\,
            I => \N__11173\
        );

    \I__2048\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__11170\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\
        );

    \I__2046\ : InMux
    port map (
            O => \N__11167\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__2045\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11161\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__11161\,
            I => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__11158\,
            I => \N__11154\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__11157\,
            I => \N__11151\
        );

    \I__2041\ : InMux
    port map (
            O => \N__11154\,
            I => \N__11146\
        );

    \I__2040\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11146\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__11146\,
            I => charx_if_generate_plus_mult1_un33_sum_i_5
        );

    \I__2038\ : InMux
    port map (
            O => \N__11143\,
            I => charx_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__2037\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11134\
        );

    \I__2036\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11134\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__11134\,
            I => un5_rowlto3_i
        );

    \I__2034\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11128\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N_575_i\
        );

    \I__2032\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11122\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__11122\,
            I => if_generate_plus_mult1_un61_sum_cry_2_s
        );

    \I__2030\ : InMux
    port map (
            O => \N__11119\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_1
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__11116\,
            I => \N__11113\
        );

    \I__2028\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11110\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__11110\,
            I => if_generate_plus_mult1_un61_sum_cry_3_s
        );

    \I__2026\ : InMux
    port map (
            O => \N__11107\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__2025\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11101\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__11101\,
            I => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\
        );

    \I__2023\ : InMux
    port map (
            O => \N__11098\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__2022\ : InMux
    port map (
            O => \N__11095\,
            I => column_1_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__2021\ : CascadeMux
    port map (
            O => \N__11092\,
            I => \N__11088\
        );

    \I__2020\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11085\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11088\,
            I => \N__11082\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__11085\,
            I => column_1_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__11082\,
            I => column_1_if_generate_plus_mult1_un54_sum_i_5
        );

    \I__2016\ : InMux
    port map (
            O => \N__11077\,
            I => charx_if_generate_plus_mult1_un33_sum_cry_1
        );

    \I__2015\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11071\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__11071\,
            I => \N_41\
        );

    \I__2013\ : CEMux
    port map (
            O => \N__11068\,
            I => \N__11062\
        );

    \I__2012\ : CEMux
    port map (
            O => \N__11067\,
            I => \N__11059\
        );

    \I__2011\ : CEMux
    port map (
            O => \N__11066\,
            I => \N__11054\
        );

    \I__2010\ : CEMux
    port map (
            O => \N__11065\,
            I => \N__11051\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__11062\,
            I => \N__11046\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__11059\,
            I => \N__11046\
        );

    \I__2007\ : CEMux
    port map (
            O => \N__11058\,
            I => \N__11043\
        );

    \I__2006\ : CEMux
    port map (
            O => \N__11057\,
            I => \N__11037\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__11054\,
            I => \N__11032\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__11051\,
            I => \N__11032\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__11046\,
            I => \N__11027\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__11043\,
            I => \N__11027\
        );

    \I__2001\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11023\
        );

    \I__2000\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11020\
        );

    \I__1999\ : InMux
    port map (
            O => \N__11040\,
            I => \N__11017\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__11037\,
            I => \N__11010\
        );

    \I__1997\ : Span4Mux_v
    port map (
            O => \N__11032\,
            I => \N__11010\
        );

    \I__1996\ : Span4Mux_s1_h
    port map (
            O => \N__11027\,
            I => \N__11010\
        );

    \I__1995\ : InMux
    port map (
            O => \N__11026\,
            I => \N__11007\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__11023\,
            I => \N__11004\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__11020\,
            I => \N__10999\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__11017\,
            I => \N__10999\
        );

    \I__1991\ : Span4Mux_h
    port map (
            O => \N__11010\,
            I => \N__10996\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__11007\,
            I => \N__10993\
        );

    \I__1989\ : Span4Mux_h
    port map (
            O => \N__11004\,
            I => \N__10990\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__10999\,
            I => \N__10985\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__10996\,
            I => \N__10985\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__10993\,
            I => un3_beamx_0
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__10990\,
            I => un3_beamx_0
        );

    \I__1984\ : Odrv4
    port map (
            O => \N__10985\,
            I => un3_beamx_0
        );

    \I__1983\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10971\
        );

    \I__1982\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10967\
        );

    \I__1981\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10964\
        );

    \I__1980\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10959\
        );

    \I__1979\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10959\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__10971\,
            I => \N__10956\
        );

    \I__1977\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10951\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10948\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__10964\,
            I => \N__10945\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__10959\,
            I => \N__10942\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__10956\,
            I => \N__10939\
        );

    \I__1972\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10934\
        );

    \I__1971\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10934\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__10951\,
            I => \N__10927\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__10948\,
            I => \N__10927\
        );

    \I__1968\ : Span4Mux_v
    port map (
            O => \N__10945\,
            I => \N__10927\
        );

    \I__1967\ : Span4Mux_s3_h
    port map (
            O => \N__10942\,
            I => \N__10924\
        );

    \I__1966\ : Sp12to4
    port map (
            O => \N__10939\,
            I => \N__10919\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10919\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__10927\,
            I => un5_beamx_0
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__10924\,
            I => un5_beamx_0
        );

    \I__1962\ : Odrv12
    port map (
            O => \N__10919\,
            I => un5_beamx_0
        );

    \I__1961\ : InMux
    port map (
            O => \N__10912\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_1
        );

    \I__1960\ : InMux
    port map (
            O => \N__10909\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__1959\ : InMux
    port map (
            O => \N__10906\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__1958\ : InMux
    port map (
            O => \N__10903\,
            I => column_1_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__10900\,
            I => \N__10897\
        );

    \I__1956\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10894\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__10894\,
            I => \column_1_if_generate_plus_mult1_un61_sum_iZ0\
        );

    \I__1954\ : InMux
    port map (
            O => \N__10891\,
            I => \N__10887\
        );

    \I__1953\ : InMux
    port map (
            O => \N__10890\,
            I => \N__10884\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__10887\,
            I => \N__10874\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__10884\,
            I => \N__10871\
        );

    \I__1950\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10860\
        );

    \I__1949\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10860\
        );

    \I__1948\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10860\
        );

    \I__1947\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10860\
        );

    \I__1946\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10860\
        );

    \I__1945\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10855\
        );

    \I__1944\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10855\
        );

    \I__1943\ : Span4Mux_s3_h
    port map (
            O => \N__10874\,
            I => \N__10852\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__10871\,
            I => \N__10847\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__10860\,
            I => \N__10847\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__10855\,
            I => \row_1_if_generate_plus_mult1_un54_sum_cZ0Z5\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__10852\,
            I => \row_1_if_generate_plus_mult1_un54_sum_cZ0Z5\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__10847\,
            I => \row_1_if_generate_plus_mult1_un54_sum_cZ0Z5\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__10840\,
            I => \un116_pixel_5_ns_1Z0Z_4_cascade_\
        );

    \I__1936\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10834\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__10834\,
            I => un116_pixel_5_ns_2
        );

    \I__1934\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10828\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__10828\,
            I => \N_362\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__10825\,
            I => \un116_pixel_7_ns_1_6_cascade_\
        );

    \I__1931\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10819\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__10819\,
            I => \N_379\
        );

    \I__1929\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10813\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__10813\,
            I => \N__10810\
        );

    \I__1927\ : Odrv12
    port map (
            O => \N__10810\,
            I => un116_pixel_3_ns_2
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__10807\,
            I => \beamY_RNI57H3N31_0Z0Z_1_cascade_\
        );

    \I__1925\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10801\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__10801\,
            I => \beamY_RNI896FQ3Z0Z_0\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__10798\,
            I => \beamY_RNI896FQ3Z0Z_0_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10792\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__10792\,
            I => \beamY_RNI57H3N31Z0Z_1\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__10789\,
            I => \un116_pixel_2_ns_1_0_6_cascade_\
        );

    \I__1919\ : InMux
    port map (
            O => \N__10786\,
            I => \N__10783\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__10783\,
            I => \beamY_RNIGO5PPVZ0Z_0\
        );

    \I__1917\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10777\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__10777\,
            I => \N_345_0_0_1\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__10774\,
            I => \font_un28_pixel_29_cascade_\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__10771\,
            I => \un116_pixel_5_am_6_cascade_\
        );

    \I__1913\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10765\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__10765\,
            I => g1_1
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__10762\,
            I => \N__10759\
        );

    \I__1910\ : InMux
    port map (
            O => \N__10759\,
            I => \N__10756\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__10756\,
            I => g0_0_x2_1
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__10753\,
            I => \un114_pixel_1_0_3__un116_pixel_2_ns_1Z0Z_2_cascade_\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__10750\,
            I => \un114_pixel_1_0_3__un116_pixel_5_ns_1Z0Z_2_cascade_\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__10747\,
            I => \N__10743\
        );

    \I__1905\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10739\
        );

    \I__1904\ : InMux
    port map (
            O => \N__10743\,
            I => \N__10736\
        );

    \I__1903\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10732\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__10739\,
            I => \N__10729\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__10736\,
            I => \N__10726\
        );

    \I__1900\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10723\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__10732\,
            I => \beamXZ0Z_9\
        );

    \I__1898\ : Odrv4
    port map (
            O => \N__10729\,
            I => \beamXZ0Z_9\
        );

    \I__1897\ : Odrv4
    port map (
            O => \N__10726\,
            I => \beamXZ0Z_9\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__10723\,
            I => \beamXZ0Z_9\
        );

    \I__1895\ : InMux
    port map (
            O => \N__10714\,
            I => un5_visiblex_cry_8
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__10711\,
            I => \un116_pixel_3_bm_2_cascade_\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__10708\,
            I => \N__10705\
        );

    \I__1892\ : InMux
    port map (
            O => \N__10705\,
            I => \N__10702\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__10702\,
            I => \un114_pixel_1_0_3__N_5_1_0\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__10699\,
            I => \un114_pixel_1_0_3__un116_pixel_4_ns_1_0_7_cascade_\
        );

    \I__1889\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10693\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__10693\,
            I => \un114_pixel_1_0_3__g2_1Z0Z_0\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__10690\,
            I => \N__10687\
        );

    \I__1886\ : InMux
    port map (
            O => \N__10687\,
            I => \N__10683\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__10686\,
            I => \N__10680\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__10683\,
            I => \N__10677\
        );

    \I__1883\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10674\
        );

    \I__1882\ : Odrv12
    port map (
            O => \N__10677\,
            I => \beamY_RNIH9THADZ0Z_4\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__10674\,
            I => \beamY_RNIH9THADZ0Z_4\
        );

    \I__1880\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10659\
        );

    \I__1879\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10655\
        );

    \I__1878\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10652\
        );

    \I__1877\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10649\
        );

    \I__1876\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10646\
        );

    \I__1875\ : InMux
    port map (
            O => \N__10664\,
            I => \N__10643\
        );

    \I__1874\ : InMux
    port map (
            O => \N__10663\,
            I => \N__10637\
        );

    \I__1873\ : InMux
    port map (
            O => \N__10662\,
            I => \N__10634\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__10659\,
            I => \N__10628\
        );

    \I__1871\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10625\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__10655\,
            I => \N__10618\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__10652\,
            I => \N__10618\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10618\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10613\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__10643\,
            I => \N__10613\
        );

    \I__1865\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10610\
        );

    \I__1864\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10605\
        );

    \I__1863\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10605\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__10637\,
            I => \N__10602\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__10634\,
            I => \N__10599\
        );

    \I__1860\ : InMux
    port map (
            O => \N__10633\,
            I => \N__10596\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__10632\,
            I => \N__10592\
        );

    \I__1858\ : InMux
    port map (
            O => \N__10631\,
            I => \N__10589\
        );

    \I__1857\ : Span12Mux_s4_v
    port map (
            O => \N__10628\,
            I => \N__10584\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10584\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__10618\,
            I => \N__10575\
        );

    \I__1854\ : Span4Mux_v
    port map (
            O => \N__10613\,
            I => \N__10575\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__10610\,
            I => \N__10575\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__10605\,
            I => \N__10575\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__10602\,
            I => \N__10568\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__10599\,
            I => \N__10568\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10568\
        );

    \I__1848\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10563\
        );

    \I__1847\ : InMux
    port map (
            O => \N__10592\,
            I => \N__10563\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__10589\,
            I => \beamYZ0Z_3\
        );

    \I__1845\ : Odrv12
    port map (
            O => \N__10584\,
            I => \beamYZ0Z_3\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__10575\,
            I => \beamYZ0Z_3\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__10568\,
            I => \beamYZ0Z_3\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__10563\,
            I => \beamYZ0Z_3\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__10552\,
            I => \N__10545\
        );

    \I__1840\ : InMux
    port map (
            O => \N__10551\,
            I => \N__10542\
        );

    \I__1839\ : InMux
    port map (
            O => \N__10550\,
            I => \N__10539\
        );

    \I__1838\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10534\
        );

    \I__1837\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10534\
        );

    \I__1836\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10531\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__10542\,
            I => \beamXZ0Z_1\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__10539\,
            I => \beamXZ0Z_1\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__10534\,
            I => \beamXZ0Z_1\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__10531\,
            I => \beamXZ0Z_1\
        );

    \I__1831\ : InMux
    port map (
            O => \N__10522\,
            I => un5_visiblex_cry_0
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__10519\,
            I => \N__10513\
        );

    \I__1829\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10510\
        );

    \I__1828\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10505\
        );

    \I__1827\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10505\
        );

    \I__1826\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10502\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__10510\,
            I => \beamXZ0Z_2\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__10505\,
            I => \beamXZ0Z_2\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__10502\,
            I => \beamXZ0Z_2\
        );

    \I__1822\ : InMux
    port map (
            O => \N__10495\,
            I => un5_visiblex_cry_1
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__10492\,
            I => \N__10487\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__10491\,
            I => \N__10482\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__10490\,
            I => \N__10479\
        );

    \I__1818\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10476\
        );

    \I__1817\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10473\
        );

    \I__1816\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10468\
        );

    \I__1815\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10468\
        );

    \I__1814\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10465\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__10476\,
            I => \beamXZ0Z_3\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__10473\,
            I => \beamXZ0Z_3\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__10468\,
            I => \beamXZ0Z_3\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__10465\,
            I => \beamXZ0Z_3\
        );

    \I__1809\ : InMux
    port map (
            O => \N__10456\,
            I => un5_visiblex_cry_2
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__10453\,
            I => \N__10445\
        );

    \I__1807\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10442\
        );

    \I__1806\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10439\
        );

    \I__1805\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10436\
        );

    \I__1804\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10431\
        );

    \I__1803\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10431\
        );

    \I__1802\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10428\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__10442\,
            I => \beamXZ0Z_4\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__10439\,
            I => \beamXZ0Z_4\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__10436\,
            I => \beamXZ0Z_4\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__10431\,
            I => \beamXZ0Z_4\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__10428\,
            I => \beamXZ0Z_4\
        );

    \I__1796\ : InMux
    port map (
            O => \N__10417\,
            I => un5_visiblex_cry_3
        );

    \I__1795\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10407\
        );

    \I__1794\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10404\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10401\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__10411\,
            I => \N__10398\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__10410\,
            I => \N__10394\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10387\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__10404\,
            I => \N__10387\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__10401\,
            I => \N__10387\
        );

    \I__1787\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10382\
        );

    \I__1786\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10382\
        );

    \I__1785\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10379\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__10387\,
            I => \beamXZ0Z_5\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__10382\,
            I => \beamXZ0Z_5\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__10379\,
            I => \beamXZ0Z_5\
        );

    \I__1781\ : InMux
    port map (
            O => \N__10372\,
            I => un5_visiblex_cry_4
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__10369\,
            I => \N__10361\
        );

    \I__1779\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10358\
        );

    \I__1778\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10355\
        );

    \I__1777\ : InMux
    port map (
            O => \N__10366\,
            I => \N__10352\
        );

    \I__1776\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10347\
        );

    \I__1775\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10347\
        );

    \I__1774\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10344\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__10358\,
            I => \beamXZ0Z_6\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__10355\,
            I => \beamXZ0Z_6\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__10352\,
            I => \beamXZ0Z_6\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__10347\,
            I => \beamXZ0Z_6\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__10344\,
            I => \beamXZ0Z_6\
        );

    \I__1768\ : InMux
    port map (
            O => \N__10333\,
            I => un5_visiblex_cry_5
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__10330\,
            I => \N__10326\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__10329\,
            I => \N__10323\
        );

    \I__1765\ : InMux
    port map (
            O => \N__10326\,
            I => \N__10316\
        );

    \I__1764\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10316\
        );

    \I__1763\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10313\
        );

    \I__1762\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10308\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__10316\,
            I => \N__10305\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__10313\,
            I => \N__10302\
        );

    \I__1759\ : InMux
    port map (
            O => \N__10312\,
            I => \N__10299\
        );

    \I__1758\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10296\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__10308\,
            I => \beamXZ0Z_7\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__10305\,
            I => \beamXZ0Z_7\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__10302\,
            I => \beamXZ0Z_7\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__10299\,
            I => \beamXZ0Z_7\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__10296\,
            I => \beamXZ0Z_7\
        );

    \I__1752\ : InMux
    port map (
            O => \N__10285\,
            I => un5_visiblex_cry_6
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__10282\,
            I => \N__10278\
        );

    \I__1750\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10274\
        );

    \I__1749\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10270\
        );

    \I__1748\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10267\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10264\
        );

    \I__1746\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10261\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__10270\,
            I => \N__10258\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__10267\,
            I => \beamXZ0Z_8\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__10264\,
            I => \beamXZ0Z_8\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10261\,
            I => \beamXZ0Z_8\
        );

    \I__1741\ : Odrv4
    port map (
            O => \N__10258\,
            I => \beamXZ0Z_8\
        );

    \I__1740\ : InMux
    port map (
            O => \N__10249\,
            I => \bfn_6_11_0_\
        );

    \I__1739\ : InMux
    port map (
            O => \N__10246\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_4
        );

    \I__1738\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10240\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__10240\,
            I => un1_beamxlt10_0
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__10237\,
            I => \N__10232\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10236\,
            I => \N__10228\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__10235\,
            I => \N__10225\
        );

    \I__1733\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10222\
        );

    \I__1732\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10219\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10216\
        );

    \I__1730\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10213\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N__10210\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__10219\,
            I => \beamXZ0Z_10\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__10216\,
            I => \beamXZ0Z_10\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__10213\,
            I => \beamXZ0Z_10\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__10210\,
            I => \beamXZ0Z_10\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__10201\,
            I => \un114_pixel_1_0_3__un3_beamxZ0Z_5_cascade_\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10195\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__10195\,
            I => \N__10192\
        );

    \I__1721\ : Odrv4
    port map (
            O => \N__10192\,
            I => \un114_pixel_1_0_3__un3_beamxZ0Z_7\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__1719\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10183\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__10183\,
            I => un18_beamylt4
        );

    \I__1717\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10176\
        );

    \I__1716\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10171\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__10176\,
            I => \N__10168\
        );

    \I__1714\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10163\
        );

    \I__1713\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10163\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__10171\,
            I => \N__10160\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__10168\,
            I => \charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__10163\,
            I => \charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__10160\,
            I => \charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__10153\,
            I => \N__10150\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10150\,
            I => \N__10147\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__10147\,
            I => \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKFZ0\
        );

    \I__1705\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10141\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__10141\,
            I => charx_if_generate_plus_mult1_un19_sum_i
        );

    \I__1703\ : InMux
    port map (
            O => \N__10138\,
            I => \N__10131\
        );

    \I__1702\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10128\
        );

    \I__1701\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10125\
        );

    \I__1700\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10120\
        );

    \I__1699\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10120\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__10131\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__10128\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__10125\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10120\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__10111\,
            I => \N__10106\
        );

    \I__1693\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10103\
        );

    \I__1692\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10098\
        );

    \I__1691\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10098\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__10103\,
            I => \beamY_RNI2MTA1Z0Z_9\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__10098\,
            I => \beamY_RNI2MTA1Z0Z_9\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__10093\,
            I => \chary_if_generate_plus_mult1_un54_sum_c4_cascade_\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10072\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10089\,
            I => \N__10072\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10088\,
            I => \N__10072\
        );

    \I__1684\ : InMux
    port map (
            O => \N__10087\,
            I => \N__10072\
        );

    \I__1683\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10065\
        );

    \I__1682\ : InMux
    port map (
            O => \N__10085\,
            I => \N__10065\
        );

    \I__1681\ : InMux
    port map (
            O => \N__10084\,
            I => \N__10065\
        );

    \I__1680\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10060\
        );

    \I__1679\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10060\
        );

    \I__1678\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10057\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__10072\,
            I => \beamY_RNICG8P9Z0Z_7\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__10065\,
            I => \beamY_RNICG8P9Z0Z_7\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__10060\,
            I => \beamY_RNICG8P9Z0Z_7\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__10057\,
            I => \beamY_RNICG8P9Z0Z_7\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10036\
        );

    \I__1672\ : InMux
    port map (
            O => \N__10047\,
            I => \N__10036\
        );

    \I__1671\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10036\
        );

    \I__1670\ : InMux
    port map (
            O => \N__10045\,
            I => \N__10031\
        );

    \I__1669\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10026\
        );

    \I__1668\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10026\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__10036\,
            I => \N__10023\
        );

    \I__1666\ : InMux
    port map (
            O => \N__10035\,
            I => \N__10018\
        );

    \I__1665\ : InMux
    port map (
            O => \N__10034\,
            I => \N__10018\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__10031\,
            I => \N__10013\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10026\,
            I => \N__10013\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__10023\,
            I => \N__10010\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__10018\,
            I => \N__10005\
        );

    \I__1660\ : Span4Mux_s2_v
    port map (
            O => \N__10013\,
            I => \N__10005\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__10010\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__10005\,
            I => chary_if_generate_plus_mult1_un61_sum_axbxc5_1
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__10000\,
            I => \un3_beamx_0_cascade_\
        );

    \I__1656\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9991\
        );

    \I__1655\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9991\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__9991\,
            I => un1_beamx_2
        );

    \I__1653\ : IoInMux
    port map (
            O => \N__9988\,
            I => \N__9985\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__9985\,
            I => \N__9982\
        );

    \I__1651\ : Span4Mux_s2_v
    port map (
            O => \N__9982\,
            I => \N__9979\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__9979\,
            I => \N__9976\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__9976\,
            I => \HSync_c\
        );

    \I__1648\ : InMux
    port map (
            O => \N__9973\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_1
        );

    \I__1647\ : InMux
    port map (
            O => \N__9970\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__9967\,
            I => \N__9964\
        );

    \I__1645\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9961\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__9961\,
            I => \N__9958\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__9958\,
            I => \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8VZ0\
        );

    \I__1642\ : InMux
    port map (
            O => \N__9955\,
            I => charx_if_generate_plus_mult1_un26_sum_cry_3
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__9952\,
            I => \N__9949\
        );

    \I__1640\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9946\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__9946\,
            I => g0_3_2
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__9943\,
            I => \beamY_RNIARUFBZ0Z_5_cascade_\
        );

    \I__1637\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9937\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__9937\,
            I => \beamY_RNIGS0LBZ0Z_5\
        );

    \I__1635\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9928\
        );

    \I__1634\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9925\
        );

    \I__1633\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9920\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__9931\,
            I => \N__9917\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__9928\,
            I => \N__9912\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__9925\,
            I => \N__9912\
        );

    \I__1629\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9903\
        );

    \I__1628\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9900\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9897\
        );

    \I__1626\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9894\
        );

    \I__1625\ : Span4Mux_h
    port map (
            O => \N__9912\,
            I => \N__9891\
        );

    \I__1624\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9882\
        );

    \I__1623\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9882\
        );

    \I__1622\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9882\
        );

    \I__1621\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9882\
        );

    \I__1620\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9877\
        );

    \I__1619\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9877\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__9903\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__9900\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__9897\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__9894\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__9891\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__9882\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__9877\,
            I => chary_if_generate_plus_mult1_un54_sum_c5
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__9862\,
            I => \chary_if_generate_plus_mult1_un54_sum_c5_cascade_\
        );

    \I__1610\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9852\
        );

    \I__1609\ : InMux
    port map (
            O => \N__9858\,
            I => \N__9847\
        );

    \I__1608\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9847\
        );

    \I__1607\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9840\
        );

    \I__1606\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9840\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__9852\,
            I => \N__9835\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__9847\,
            I => \N__9835\
        );

    \I__1603\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9830\
        );

    \I__1602\ : InMux
    port map (
            O => \N__9845\,
            I => \N__9830\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__9840\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__9835\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__9830\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0
        );

    \I__1598\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9820\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__9820\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0_0
        );

    \I__1596\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9812\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__9816\,
            I => \N__9809\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__9815\,
            I => \N__9805\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__9812\,
            I => \N__9800\
        );

    \I__1592\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9789\
        );

    \I__1591\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9789\
        );

    \I__1590\ : InMux
    port map (
            O => \N__9805\,
            I => \N__9789\
        );

    \I__1589\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9789\
        );

    \I__1588\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9789\
        );

    \I__1587\ : Odrv4
    port map (
            O => \N__9800\,
            I => \beamY_RNIDO3IZ0Z_9\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__9789\,
            I => \beamY_RNIDO3IZ0Z_9\
        );

    \I__1585\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9777\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__9783\,
            I => \N__9774\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__9782\,
            I => \N__9771\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__9781\,
            I => \N__9766\
        );

    \I__1581\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9757\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__9777\,
            I => \N__9754\
        );

    \I__1579\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9751\
        );

    \I__1578\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9746\
        );

    \I__1577\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9746\
        );

    \I__1576\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9743\
        );

    \I__1575\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9740\
        );

    \I__1574\ : InMux
    port map (
            O => \N__9765\,
            I => \N__9735\
        );

    \I__1573\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9730\
        );

    \I__1572\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9730\
        );

    \I__1571\ : InMux
    port map (
            O => \N__9762\,
            I => \N__9725\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9725\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__9760\,
            I => \N__9722\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__9757\,
            I => \N__9715\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__9754\,
            I => \N__9715\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9706\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__9746\,
            I => \N__9706\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__9743\,
            I => \N__9706\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__9740\,
            I => \N__9706\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__9739\,
            I => \N__9703\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__9738\,
            I => \N__9700\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__9735\,
            I => \N__9695\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__9730\,
            I => \N__9690\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__9725\,
            I => \N__9690\
        );

    \I__1557\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9685\
        );

    \I__1556\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9685\
        );

    \I__1555\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9682\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__9715\,
            I => \N__9677\
        );

    \I__1553\ : Span4Mux_v
    port map (
            O => \N__9706\,
            I => \N__9677\
        );

    \I__1552\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9672\
        );

    \I__1551\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9672\
        );

    \I__1550\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9669\
        );

    \I__1549\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9666\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__9695\,
            I => \N__9661\
        );

    \I__1547\ : Span4Mux_v
    port map (
            O => \N__9690\,
            I => \N__9661\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__9685\,
            I => \N__9652\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__9682\,
            I => \N__9652\
        );

    \I__1544\ : Sp12to4
    port map (
            O => \N__9677\,
            I => \N__9652\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__9672\,
            I => \N__9652\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__9669\,
            I => \N__9647\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__9666\,
            I => \N__9647\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__9661\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1539\ : Odrv12
    port map (
            O => \N__9652\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1538\ : Odrv12
    port map (
            O => \N__9647\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__9640\,
            I => \N__9635\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__9639\,
            I => \N__9631\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__9638\,
            I => \N__9627\
        );

    \I__1534\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9621\
        );

    \I__1533\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9621\
        );

    \I__1532\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9618\
        );

    \I__1531\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9611\
        );

    \I__1530\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9611\
        );

    \I__1529\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9611\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__9621\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__9618\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__9611\,
            I => chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__9604\,
            I => \N__9601\
        );

    \I__1524\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9598\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__9598\,
            I => \N__9595\
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__9595\,
            I => g0_4_2
        );

    \I__1521\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9584\
        );

    \I__1520\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9579\
        );

    \I__1519\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9579\
        );

    \I__1518\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9572\
        );

    \I__1517\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9572\
        );

    \I__1516\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9572\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__9584\,
            I => \N__9565\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__9579\,
            I => \N__9565\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9562\
        );

    \I__1512\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9559\
        );

    \I__1511\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9556\
        );

    \I__1510\ : Span4Mux_v
    port map (
            O => \N__9565\,
            I => \N__9551\
        );

    \I__1509\ : Span4Mux_h
    port map (
            O => \N__9562\,
            I => \N__9551\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__9559\,
            I => \N__9546\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__9556\,
            I => \N__9546\
        );

    \I__1506\ : Span4Mux_h
    port map (
            O => \N__9551\,
            I => \N__9530\
        );

    \I__1505\ : Span4Mux_h
    port map (
            O => \N__9546\,
            I => \N__9530\
        );

    \I__1504\ : InMux
    port map (
            O => \N__9545\,
            I => \N__9521\
        );

    \I__1503\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9521\
        );

    \I__1502\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9521\
        );

    \I__1501\ : InMux
    port map (
            O => \N__9542\,
            I => \N__9521\
        );

    \I__1500\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9512\
        );

    \I__1499\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9512\
        );

    \I__1498\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9512\
        );

    \I__1497\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9512\
        );

    \I__1496\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9507\
        );

    \I__1495\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9507\
        );

    \I__1494\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9504\
        );

    \I__1493\ : Span4Mux_v
    port map (
            O => \N__9530\,
            I => \N__9501\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__9521\,
            I => \N__9496\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__9512\,
            I => \N__9496\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9491\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__9504\,
            I => \N__9491\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__9501\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1487\ : Odrv12
    port map (
            O => \N__9496\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1486\ : Odrv12
    port map (
            O => \N__9491\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__9484\,
            I => \N__9481\
        );

    \I__1484\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9475\
        );

    \I__1483\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9468\
        );

    \I__1482\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9468\
        );

    \I__1481\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9468\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__9475\,
            I => chary_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__9468\,
            I => chary_if_generate_plus_mult1_un54_sum_axb3
        );

    \I__1478\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9455\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__9462\,
            I => \N__9452\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__9461\,
            I => \N__9442\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__9460\,
            I => \N__9439\
        );

    \I__1474\ : InMux
    port map (
            O => \N__9459\,
            I => \N__9434\
        );

    \I__1473\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9434\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9431\
        );

    \I__1471\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9428\
        );

    \I__1470\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9422\
        );

    \I__1469\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9422\
        );

    \I__1468\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9413\
        );

    \I__1467\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9413\
        );

    \I__1466\ : InMux
    port map (
            O => \N__9447\,
            I => \N__9413\
        );

    \I__1465\ : InMux
    port map (
            O => \N__9446\,
            I => \N__9413\
        );

    \I__1464\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9408\
        );

    \I__1463\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9408\
        );

    \I__1462\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9405\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9400\
        );

    \I__1460\ : Span4Mux_v
    port map (
            O => \N__9431\,
            I => \N__9395\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__9428\,
            I => \N__9395\
        );

    \I__1458\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9392\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__9422\,
            I => \N__9389\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__9413\,
            I => \N__9382\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__9408\,
            I => \N__9382\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9382\
        );

    \I__1453\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9377\
        );

    \I__1452\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9377\
        );

    \I__1451\ : Span4Mux_v
    port map (
            O => \N__9400\,
            I => \N__9372\
        );

    \I__1450\ : Span4Mux_v
    port map (
            O => \N__9395\,
            I => \N__9372\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__9392\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__9389\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1447\ : Odrv12
    port map (
            O => \N__9382\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__9377\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__9372\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum
        );

    \I__1444\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9354\
        );

    \I__1443\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9349\
        );

    \I__1442\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9349\
        );

    \I__1441\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9345\
        );

    \I__1440\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9342\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__9354\,
            I => \N__9337\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__9349\,
            I => \N__9337\
        );

    \I__1437\ : InMux
    port map (
            O => \N__9348\,
            I => \N__9334\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__9345\,
            I => \beamY_RNITFRN03Z0Z_5\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__9342\,
            I => \beamY_RNITFRN03Z0Z_5\
        );

    \I__1434\ : Odrv4
    port map (
            O => \N__9337\,
            I => \beamY_RNITFRN03Z0Z_5\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__9334\,
            I => \beamY_RNITFRN03Z0Z_5\
        );

    \I__1432\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9319\
        );

    \I__1431\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9314\
        );

    \I__1430\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9314\
        );

    \I__1429\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9311\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N__9308\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__9314\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__9311\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__9308\,
            I => chary_if_generate_plus_mult1_un75_sum_c5
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__9301\,
            I => \beamY_RNIH9THADZ0Z_4_cascade_\
        );

    \I__1423\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9292\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__9297\,
            I => \N__9289\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9286\
        );

    \I__1420\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9283\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__9292\,
            I => \N__9279\
        );

    \I__1418\ : InMux
    port map (
            O => \N__9289\,
            I => \N__9276\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__9286\,
            I => \N__9271\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__9283\,
            I => \N__9271\
        );

    \I__1415\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9268\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__9279\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__9276\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0
        );

    \I__1412\ : Odrv4
    port map (
            O => \N__9271\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__9268\,
            I => chary_if_generate_plus_mult1_un61_sum_axb3_0
        );

    \I__1410\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9251\
        );

    \I__1409\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9248\
        );

    \I__1408\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9245\
        );

    \I__1407\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9240\
        );

    \I__1406\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9240\
        );

    \I__1405\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9237\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__9251\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_d
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__9248\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_d
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__9245\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_d
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__9240\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_d
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__9237\,
            I => chary_if_generate_plus_mult1_un61_sum_ac0_7_d
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__1398\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9216\
        );

    \I__1397\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9216\
        );

    \I__1396\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9213\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__9216\,
            I => \N__9210\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__9213\,
            I => \N__9207\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__9210\,
            I => \N__9204\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__9207\,
            I => \beamY_RNIKHPCA1Z0Z_4\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__9204\,
            I => \beamY_RNIKHPCA1Z0Z_4\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__9199\,
            I => \chary_if_generate_plus_mult1_un61_sum_ac0_7_d_cascade_\
        );

    \I__1389\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9193\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__9193\,
            I => chary_if_generate_plus_mult1_un68_sum_axb4
        );

    \I__1387\ : InMux
    port map (
            O => \N__9190\,
            I => \N__9187\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__9187\,
            I => \N__9181\
        );

    \I__1385\ : InMux
    port map (
            O => \N__9186\,
            I => \N__9178\
        );

    \I__1384\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9173\
        );

    \I__1383\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9173\
        );

    \I__1382\ : Span4Mux_v
    port map (
            O => \N__9181\,
            I => \N__9170\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__9178\,
            I => \beamY_RNI2TEJF4Z0Z_4\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__9173\,
            I => \beamY_RNI2TEJF4Z0Z_4\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__9170\,
            I => \beamY_RNI2TEJF4Z0Z_4\
        );

    \I__1378\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9154\
        );

    \I__1377\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9154\
        );

    \I__1376\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9151\
        );

    \I__1375\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9146\
        );

    \I__1374\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9146\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__9154\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__9151\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__9146\,
            I => chary_if_generate_plus_mult1_un68_sum_c4
        );

    \I__1370\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9134\
        );

    \I__1369\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9131\
        );

    \I__1368\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9128\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__9134\,
            I => \N__9125\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__9131\,
            I => chary_if_generate_plus_mult1_un61_sum_axb4_0
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__9128\,
            I => chary_if_generate_plus_mult1_un61_sum_axb4_0
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__9125\,
            I => chary_if_generate_plus_mult1_un61_sum_axb4_0
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__9118\,
            I => \g0_0_x2_1_1_cascade_\
        );

    \I__1362\ : CascadeMux
    port map (
            O => \N__9115\,
            I => \beamY_RNI2TEJF4Z0Z_4_cascade_\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__9112\,
            I => \N__9109\
        );

    \I__1360\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__9106\,
            I => \un114_pixel_1_0_3__g0_8Z0Z_1\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__9103\,
            I => \chary_if_generate_plus_mult1_un61_sum_0_3_cascade_\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__9100\,
            I => \un114_pixel_1_0_3__g0_1Z0Z_1_cascade_\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9094\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__9094\,
            I => chary_if_generate_plus_mult1_un61_sum_0_3
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__9091\,
            I => \un114_pixel_1_0_3__g0_3Z0Z_0_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9085\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__9085\,
            I => chary_if_generate_plus_mult1_un75_sum_i_0_5
        );

    \I__1351\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9078\
        );

    \I__1350\ : InMux
    port map (
            O => \N__9081\,
            I => \N__9075\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__9078\,
            I => chary_if_generate_plus_mult1_un68_sum_c4_0
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__9075\,
            I => chary_if_generate_plus_mult1_un68_sum_c4_0
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__9070\,
            I => \un114_pixel_1_0_3__g0Z0Z_1_cascade_\
        );

    \I__1346\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9064\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__9064\,
            I => chary_if_generate_plus_mult1_un68_sum_0_0_0_0_5
        );

    \I__1344\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9058\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__9058\,
            I => g2
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__9055\,
            I => \un114_pixel_1_0_3__g0Z0Z_3_cascade_\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__1340\ : InMux
    port map (
            O => \N__9049\,
            I => \N__9046\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__9046\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__9043\,
            I => \N__9040\
        );

    \I__1337\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9037\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__9037\,
            I => \N__9034\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__9034\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i
        );

    \I__1334\ : InMux
    port map (
            O => \N__9031\,
            I => \N__9028\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__9028\,
            I => counter_27
        );

    \I__1332\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9016\
        );

    \I__1331\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9016\
        );

    \I__1330\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9013\
        );

    \I__1329\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9008\
        );

    \I__1328\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9008\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__9016\,
            I => \counterZ0Z_5\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__9013\,
            I => \counterZ0Z_5\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__9008\,
            I => \counterZ0Z_5\
        );

    \I__1324\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8995\
        );

    \I__1323\ : InMux
    port map (
            O => \N__9000\,
            I => \N__8995\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__8995\,
            I => slaveselect_1_0_4
        );

    \I__1321\ : IoInMux
    port map (
            O => \N__8992\,
            I => \N__8988\
        );

    \I__1320\ : IoInMux
    port map (
            O => \N__8991\,
            I => \N__8985\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8980\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8980\
        );

    \I__1317\ : IoSpan4Mux
    port map (
            O => \N__8980\,
            I => \N__8977\
        );

    \I__1316\ : Span4Mux_s3_v
    port map (
            O => \N__8977\,
            I => \N__8974\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__8974\,
            I => un1_slaveselect_1_i
        );

    \I__1314\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8959\
        );

    \I__1313\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8959\
        );

    \I__1312\ : InMux
    port map (
            O => \N__8969\,
            I => \N__8959\
        );

    \I__1311\ : InMux
    port map (
            O => \N__8968\,
            I => \N__8952\
        );

    \I__1310\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8952\
        );

    \I__1309\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8952\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__8959\,
            I => un3_slaveselect
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__8952\,
            I => un3_slaveselect
        );

    \I__1306\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8944\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__8944\,
            I => counter_28
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__8941\,
            I => \N__8934\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__8940\,
            I => \N__8931\
        );

    \I__1302\ : InMux
    port map (
            O => \N__8939\,
            I => \N__8928\
        );

    \I__1301\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8923\
        );

    \I__1300\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8923\
        );

    \I__1299\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8918\
        );

    \I__1298\ : InMux
    port map (
            O => \N__8931\,
            I => \N__8918\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__8928\,
            I => \counterZ0Z_4\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__8923\,
            I => \counterZ0Z_4\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__8918\,
            I => \counterZ0Z_4\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__8911\,
            I => \N__8904\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__8910\,
            I => \N__8901\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__8909\,
            I => \N__8895\
        );

    \I__1291\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8890\
        );

    \I__1290\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8883\
        );

    \I__1289\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8883\
        );

    \I__1288\ : InMux
    port map (
            O => \N__8901\,
            I => \N__8883\
        );

    \I__1287\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8880\
        );

    \I__1286\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8869\
        );

    \I__1285\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8869\
        );

    \I__1284\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8869\
        );

    \I__1283\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8869\
        );

    \I__1282\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8869\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__8890\,
            I => \slaveselectZ0\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__8883\,
            I => \slaveselectZ0\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__8880\,
            I => \slaveselectZ0\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__8869\,
            I => \slaveselectZ0\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__8860\,
            I => \N__8855\
        );

    \I__1276\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8847\
        );

    \I__1275\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8844\
        );

    \I__1274\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8839\
        );

    \I__1273\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8839\
        );

    \I__1272\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8836\
        );

    \I__1271\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8829\
        );

    \I__1270\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8829\
        );

    \I__1269\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8829\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__8847\,
            I => un1_counter_0
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__8844\,
            I => un1_counter_0
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__8839\,
            I => un1_counter_0
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__8836\,
            I => un1_counter_0
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__8829\,
            I => un1_counter_0
        );

    \I__1263\ : IoInMux
    port map (
            O => \N__8818\,
            I => \N__8814\
        );

    \I__1262\ : IoInMux
    port map (
            O => \N__8817\,
            I => \N__8811\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__8814\,
            I => \N__8806\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8806\
        );

    \I__1259\ : Span4Mux_s2_v
    port map (
            O => \N__8806\,
            I => \N__8803\
        );

    \I__1258\ : Sp12to4
    port map (
            O => \N__8803\,
            I => \N__8799\
        );

    \I__1257\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8796\
        );

    \I__1256\ : Odrv12
    port map (
            O => \N__8799\,
            I => \nCS1_c\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__8796\,
            I => \nCS1_c\
        );

    \I__1254\ : SRMux
    port map (
            O => \N__8791\,
            I => \N__8788\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__8788\,
            I => \N__8785\
        );

    \I__1252\ : Span4Mux_h
    port map (
            O => \N__8785\,
            I => \N__8782\
        );

    \I__1251\ : Odrv4
    port map (
            O => \N__8782\,
            I => \nCS1_0_sqmuxa\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8779\,
            I => un8_beamx_cry_6
        );

    \I__1249\ : InMux
    port map (
            O => \N__8776\,
            I => un8_beamx_cry_7
        );

    \I__1248\ : InMux
    port map (
            O => \N__8773\,
            I => \bfn_5_10_0_\
        );

    \I__1247\ : InMux
    port map (
            O => \N__8770\,
            I => un8_beamx_cry_9
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__8767\,
            I => \N__8764\
        );

    \I__1245\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8761\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__8761\,
            I => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0\
        );

    \I__1243\ : InMux
    port map (
            O => \N__8758\,
            I => charx_if_generate_plus_mult1_un19_sum_cry_2
        );

    \I__1242\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8752\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__8752\,
            I => un13_beamylt7
        );

    \I__1240\ : CascadeMux
    port map (
            O => \N__8749\,
            I => \N__8745\
        );

    \I__1239\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8740\
        );

    \I__1238\ : InMux
    port map (
            O => \N__8745\,
            I => \N__8740\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__8740\,
            I => if_generate_plus_mult1_un75_sum_axbxc5
        );

    \I__1236\ : InMux
    port map (
            O => \N__8737\,
            I => \N__8733\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8730\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__8733\,
            I => if_generate_plus_mult1_un75_sum_axbxc3
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__8730\,
            I => if_generate_plus_mult1_un75_sum_axbxc3
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__8725\,
            I => \row_1_if_generate_plus_mult1_un82_sum_axb4_i_cascade_\
        );

    \I__1231\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8719\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__8719\,
            I => \row_1_if_generate_plus_mult1_un82_sum_ac0_7_0Z0Z_1\
        );

    \I__1229\ : InMux
    port map (
            O => \N__8716\,
            I => un8_beamx_cry_1
        );

    \I__1228\ : InMux
    port map (
            O => \N__8713\,
            I => un8_beamx_cry_2
        );

    \I__1227\ : InMux
    port map (
            O => \N__8710\,
            I => un8_beamx_cry_3
        );

    \I__1226\ : InMux
    port map (
            O => \N__8707\,
            I => un8_beamx_cry_4
        );

    \I__1225\ : InMux
    port map (
            O => \N__8704\,
            I => un8_beamx_cry_5
        );

    \I__1224\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8692\
        );

    \I__1223\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8692\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8692\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__8692\,
            I => chary_if_generate_plus_mult1_un47_sum_c5
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__8689\,
            I => \beamY_RNITURI3_0Z0Z_7_cascade_\
        );

    \I__1219\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8683\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__8683\,
            I => \beamY_RNITURI3Z0Z_7\
        );

    \I__1217\ : InMux
    port map (
            O => \N__8680\,
            I => \N__8677\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__8677\,
            I => un4_beamy_0
        );

    \I__1215\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8671\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__8671\,
            I => un8_beamy
        );

    \I__1213\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8665\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__8665\,
            I => \un114_pixel_1_0_3__un15_beamyZ0Z_2\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__8662\,
            I => \un1_beamx_2_cascade_\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__8659\,
            I => \N__8656\
        );

    \I__1209\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8653\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__8653\,
            I => \N__8650\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__8650\,
            I => \un114_pixel_1_0_3__un5_beamxZ0Z_3\
        );

    \I__1206\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8638\
        );

    \I__1205\ : InMux
    port map (
            O => \N__8646\,
            I => \N__8635\
        );

    \I__1204\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8630\
        );

    \I__1203\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8630\
        );

    \I__1202\ : InMux
    port map (
            O => \N__8643\,
            I => \N__8626\
        );

    \I__1201\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8621\
        );

    \I__1200\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8621\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__8638\,
            I => \N__8617\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__8635\,
            I => \N__8612\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__8630\,
            I => \N__8612\
        );

    \I__1196\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8609\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__8626\,
            I => \N__8602\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__8621\,
            I => \N__8602\
        );

    \I__1193\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8596\
        );

    \I__1192\ : Span4Mux_v
    port map (
            O => \N__8617\,
            I => \N__8589\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__8612\,
            I => \N__8589\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8589\
        );

    \I__1189\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8584\
        );

    \I__1188\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8584\
        );

    \I__1187\ : Span4Mux_h
    port map (
            O => \N__8602\,
            I => \N__8581\
        );

    \I__1186\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8574\
        );

    \I__1185\ : InMux
    port map (
            O => \N__8600\,
            I => \N__8574\
        );

    \I__1184\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8574\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__8596\,
            I => \beamYZ0Z_4\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__8589\,
            I => \beamYZ0Z_4\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__8584\,
            I => \beamYZ0Z_4\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__8581\,
            I => \beamYZ0Z_4\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__8574\,
            I => \beamYZ0Z_4\
        );

    \I__1178\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8560\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__8560\,
            I => \un114_pixel_1_0_3__g0_1Z0Z_3\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__8557\,
            I => \un114_pixel_1_0_3__un18_beamylto9Z0Z_2_cascade_\
        );

    \I__1175\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__8551\,
            I => un18_beamylt10_0
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__8548\,
            I => \N__8542\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__8547\,
            I => \N__8539\
        );

    \I__1171\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8536\
        );

    \I__1170\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8533\
        );

    \I__1169\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8530\
        );

    \I__1168\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8527\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__8536\,
            I => \N__8524\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__8533\,
            I => \N__8515\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__8530\,
            I => \N__8515\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__8527\,
            I => \N__8515\
        );

    \I__1163\ : Span4Mux_h
    port map (
            O => \N__8524\,
            I => \N__8512\
        );

    \I__1162\ : InMux
    port map (
            O => \N__8523\,
            I => \N__8509\
        );

    \I__1161\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8506\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__8515\,
            I => \N__8501\
        );

    \I__1159\ : Span4Mux_v
    port map (
            O => \N__8512\,
            I => \N__8501\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8498\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8495\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__8501\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__8498\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1154\ : Odrv12
    port map (
            O => \N__8495\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__8488\,
            I => \beamY_RNINITP61Z0Z_5_cascade_\
        );

    \I__1152\ : InMux
    port map (
            O => \N__8485\,
            I => \N__8482\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__8482\,
            I => \beamY_RNINITP61_1Z0Z_5\
        );

    \I__1150\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8473\
        );

    \I__1149\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8473\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__8473\,
            I => chary_if_generate_plus_mult1_un40_sum_axb3
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__8470\,
            I => \chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0_cascade_\
        );

    \I__1146\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8464\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__8464\,
            I => chary_if_generate_plus_mult1_un47_sum_axbxc5_2
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__8461\,
            I => \chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_\
        );

    \I__1143\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8446\
        );

    \I__1142\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8446\
        );

    \I__1141\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8446\
        );

    \I__1140\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8446\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__8446\,
            I => chary_if_generate_plus_mult1_un40_sum_c4
        );

    \I__1138\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8440\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__8440\,
            I => un5_visibley_0_29
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__8437\,
            I => \chary_if_generate_plus_mult1_un61_sum_c5_cascade_\
        );

    \I__1135\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8428\
        );

    \I__1134\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8428\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__8428\,
            I => chary_if_generate_plus_mult1_un61_sum_0_1_5
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__8425\,
            I => \chary_if_generate_plus_mult1_un68_sum_c4_0_cascade_\
        );

    \I__1131\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8419\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__8419\,
            I => g0_0_3
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__8416\,
            I => \g1_0_cascade_\
        );

    \I__1128\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8410\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8407\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__8407\,
            I => un4_beamylt6
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__8404\,
            I => \chary_if_generate_plus_mult1_un75_sum_c5_N_9_cascade_\
        );

    \I__1124\ : InMux
    port map (
            O => \N__8401\,
            I => \N__8398\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__8398\,
            I => g0_1_2
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__8395\,
            I => \N__8392\
        );

    \I__1121\ : InMux
    port map (
            O => \N__8392\,
            I => \N__8389\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__8389\,
            I => \N__8386\
        );

    \I__1119\ : Span4Mux_h
    port map (
            O => \N__8386\,
            I => \N__8383\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__8380\,
            I => g0_2_0
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__8377\,
            I => \N__8374\
        );

    \I__1115\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__8371\,
            I => chary_if_generate_plus_mult1_un61_sum_1_0_1_0_3
        );

    \I__1113\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8363\
        );

    \I__1112\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8360\
        );

    \I__1111\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8357\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__8363\,
            I => \counterZ0Z_3\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__8360\,
            I => \counterZ0Z_3\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__8357\,
            I => \counterZ0Z_3\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__8350\,
            I => \N__8344\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__8349\,
            I => \N__8341\
        );

    \I__1105\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8336\
        );

    \I__1104\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8336\
        );

    \I__1103\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8333\
        );

    \I__1102\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8330\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__8336\,
            I => \counterZ0Z_1\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__8333\,
            I => \counterZ0Z_1\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__8330\,
            I => \counterZ0Z_1\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__8323\,
            I => \un1_counterlto3_0_cascade_\
        );

    \I__1097\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8313\
        );

    \I__1096\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8313\
        );

    \I__1095\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8310\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__8313\,
            I => \N__8307\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__8310\,
            I => \counterZ0Z_2\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__8307\,
            I => \counterZ0Z_2\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__8302\,
            I => \g0_0_1_cascade_\
        );

    \I__1090\ : InMux
    port map (
            O => \N__8299\,
            I => \N__8296\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__8296\,
            I => chary_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1088\ : InMux
    port map (
            O => \N__8293\,
            I => counter_cry_3
        );

    \I__1087\ : InMux
    port map (
            O => \N__8290\,
            I => counter_cry_4
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__8287\,
            I => \slaveselect_1_0_4_cascade_\
        );

    \I__1085\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__8281\,
            I => counter_30
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__8278\,
            I => \un3_slaveselect_cascade_\
        );

    \I__1082\ : InMux
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__8272\,
            I => counter_29
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__8269\,
            I => \counter_31_cascade_\
        );

    \I__1079\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8258\
        );

    \I__1078\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8258\
        );

    \I__1077\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8253\
        );

    \I__1076\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8253\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__8258\,
            I => \counterZ0Z_0\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__8253\,
            I => \counterZ0Z_0\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__8248\,
            I => \N__8245\
        );

    \I__1072\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8242\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8239\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__8239\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KCZ0Z4\
        );

    \I__1069\ : InMux
    port map (
            O => \N__8236\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__8233\,
            I => \N__8230\
        );

    \I__1067\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8227\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__8227\,
            I => \N__8224\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__8224\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGSZ0Z6\
        );

    \I__1064\ : InMux
    port map (
            O => \N__8221\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__1063\ : InMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8212\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__8212\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8
        );

    \I__1060\ : InMux
    port map (
            O => \N__8209\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__1059\ : InMux
    port map (
            O => \N__8206\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7
        );

    \I__1058\ : InMux
    port map (
            O => \N__8203\,
            I => \N__8196\
        );

    \I__1057\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8196\
        );

    \I__1056\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8193\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__8196\,
            I => \N__8190\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__8193\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__8190\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7\
        );

    \I__1052\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8179\
        );

    \I__1051\ : InMux
    port map (
            O => \N__8184\,
            I => \N__8179\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__8179\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8
        );

    \I__1049\ : InMux
    port map (
            O => \N__8176\,
            I => counter_cry_1
        );

    \I__1048\ : InMux
    port map (
            O => \N__8173\,
            I => counter_cry_2
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__8170\,
            I => \N__8167\
        );

    \I__1046\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__1044\ : Odrv12
    port map (
            O => \N__8161\,
            I => \row_1_if_generate_plus_mult1_un68_sum_c5_0_nsZ0Z_1\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__8158\,
            I => \N__8154\
        );

    \I__1042\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8149\
        );

    \I__1041\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8144\
        );

    \I__1040\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8144\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8141\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__8149\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__8144\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__8141\,
            I => row_1_if_generate_plus_mult1_un68_sum_c5
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__8134\,
            I => \row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0_cascade_\
        );

    \I__1034\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8128\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__8128\,
            I => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5\
        );

    \I__1032\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8121\
        );

    \I__1031\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8118\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__8121\,
            I => if_generate_plus_mult1_un54_sum_axbxc3
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__8118\,
            I => if_generate_plus_mult1_un54_sum_axbxc3
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__8113\,
            I => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5_cascade_\
        );

    \I__1027\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8107\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__8107\,
            I => row_1_if_generate_plus_mult1_un61_sum_c5
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__8104\,
            I => \row_1_if_generate_plus_mult1_un61_sum_c5_cascade_\
        );

    \I__1024\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8098\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__8098\,
            I => \row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__8092\,
            I => if_generate_plus_mult1_un68_sum_c5_0_bm
        );

    \I__1020\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8086\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__8086\,
            I => \N__8083\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__8083\,
            I => row_1_if_generate_plus_mult1_un61_sum_ac0_7_c
        );

    \I__1017\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8074\
        );

    \I__1016\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8074\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__8074\,
            I => \row_1_if_generate_plus_mult1_un75_sum_cZ0Z4\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__8071\,
            I => \row_1_if_generate_plus_mult1_un75_sum_cZ0Z4_cascade_\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__8068\,
            I => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_\
        );

    \I__1012\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8056\
        );

    \I__1011\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8056\
        );

    \I__1010\ : InMux
    port map (
            O => \N__8063\,
            I => \N__8056\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__8056\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__8053\,
            I => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_\
        );

    \I__1007\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8041\
        );

    \I__1006\ : InMux
    port map (
            O => \N__8049\,
            I => \N__8041\
        );

    \I__1005\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8041\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8041\,
            I => if_generate_plus_mult1_un68_sum_axbxc3
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__8038\,
            I => \N__8035\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8035\,
            I => \N__8032\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__8032\,
            I => un5_visibley_c5
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__8029\,
            I => \un5_visibley_c5_cascade_\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__8026\,
            I => \un114_pixel_1_0_3__un5_beamxZ0Z_5_cascade_\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__8023\,
            I => \un114_pixel_1_0_3__g0_1Z0Z_0_cascade_\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__8020\,
            I => \N__8017\
        );

    \I__996\ : InMux
    port map (
            O => \N__8017\,
            I => \N__8014\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__8014\,
            I => \N__8011\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__8011\,
            I => un4_beamylt8_0
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__8008\,
            I => \N__8005\
        );

    \I__992\ : InMux
    port map (
            O => \N__8005\,
            I => \N__8001\
        );

    \I__991\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7998\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__8001\,
            I => \N__7995\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7991\
        );

    \I__988\ : Span4Mux_h
    port map (
            O => \N__7995\,
            I => \N__7988\
        );

    \I__987\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7985\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__7991\,
            I => un5_visibley_c2
        );

    \I__985\ : Odrv4
    port map (
            O => \N__7988\,
            I => un5_visibley_c2
        );

    \I__984\ : LocalMux
    port map (
            O => \N__7985\,
            I => un5_visibley_c2
        );

    \I__983\ : InMux
    port map (
            O => \N__7978\,
            I => \N__7972\
        );

    \I__982\ : InMux
    port map (
            O => \N__7977\,
            I => \N__7969\
        );

    \I__981\ : InMux
    port map (
            O => \N__7976\,
            I => \N__7964\
        );

    \I__980\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7964\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__7972\,
            I => \N__7961\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__7969\,
            I => \N__7956\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__7964\,
            I => \N__7956\
        );

    \I__976\ : Span4Mux_h
    port map (
            O => \N__7961\,
            I => \N__7952\
        );

    \I__975\ : Span4Mux_h
    port map (
            O => \N__7956\,
            I => \N__7949\
        );

    \I__974\ : InMux
    port map (
            O => \N__7955\,
            I => \N__7946\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__7952\,
            I => un1_beamy_4
        );

    \I__972\ : Odrv4
    port map (
            O => \N__7949\,
            I => un1_beamy_4
        );

    \I__971\ : LocalMux
    port map (
            O => \N__7946\,
            I => un1_beamy_4
        );

    \I__970\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7933\
        );

    \I__969\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7926\
        );

    \I__968\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7926\
        );

    \I__967\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7926\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__7933\,
            I => \N__7917\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__7926\,
            I => \N__7917\
        );

    \I__964\ : InMux
    port map (
            O => \N__7925\,
            I => \N__7912\
        );

    \I__963\ : InMux
    port map (
            O => \N__7924\,
            I => \N__7912\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7907\
        );

    \I__961\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7903\
        );

    \I__960\ : Span4Mux_h
    port map (
            O => \N__7917\,
            I => \N__7900\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__7912\,
            I => \N__7897\
        );

    \I__958\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7894\
        );

    \I__957\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7887\
        );

    \I__956\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7887\
        );

    \I__955\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7887\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__7903\,
            I => \beamYZ0Z_8\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__7900\,
            I => \beamYZ0Z_8\
        );

    \I__952\ : Odrv12
    port map (
            O => \N__7897\,
            I => \beamYZ0Z_8\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__7894\,
            I => \beamYZ0Z_8\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__7887\,
            I => \beamYZ0Z_8\
        );

    \I__949\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7867\
        );

    \I__948\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7860\
        );

    \I__947\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7860\
        );

    \I__946\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7860\
        );

    \I__945\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7853\
        );

    \I__944\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7853\
        );

    \I__943\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7853\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__7867\,
            I => \N__7845\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__7860\,
            I => \N__7845\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__7853\,
            I => \N__7845\
        );

    \I__939\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7841\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__7845\,
            I => \N__7838\
        );

    \I__937\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7835\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__7841\,
            I => \beamYZ0Z_9\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__7838\,
            I => \beamYZ0Z_9\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__7835\,
            I => \beamYZ0Z_9\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__7828\,
            I => \un114_pixel_1_0_3__un8_beamylto9Z0Z_1_cascade_\
        );

    \I__932\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7820\
        );

    \I__931\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7811\
        );

    \I__930\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7811\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7806\
        );

    \I__928\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7797\
        );

    \I__927\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7797\
        );

    \I__926\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7797\
        );

    \I__925\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7797\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__7811\,
            I => \N__7794\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__7810\,
            I => \N__7791\
        );

    \I__922\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7788\
        );

    \I__921\ : Span4Mux_v
    port map (
            O => \N__7806\,
            I => \N__7783\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__7797\,
            I => \N__7783\
        );

    \I__919\ : Span4Mux_h
    port map (
            O => \N__7794\,
            I => \N__7780\
        );

    \I__918\ : InMux
    port map (
            O => \N__7791\,
            I => \N__7777\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__7788\,
            I => \beamYZ0Z_7\
        );

    \I__916\ : Odrv4
    port map (
            O => \N__7783\,
            I => \beamYZ0Z_7\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__7780\,
            I => \beamYZ0Z_7\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7777\,
            I => \beamYZ0Z_7\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__7768\,
            I => \un114_pixel_1_0_3__un1_beamylto9Z0Z_0_cascade_\
        );

    \I__912\ : CascadeMux
    port map (
            O => \N__7765\,
            I => \un4_beamylt6_cascade_\
        );

    \I__911\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7759\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__7759\,
            I => \N__7755\
        );

    \I__909\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7752\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__7755\,
            I => un5_visibley_ac0_11_d
        );

    \I__907\ : LocalMux
    port map (
            O => \N__7752\,
            I => un5_visibley_ac0_11_d
        );

    \I__906\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7744\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__7744\,
            I => \N__7740\
        );

    \I__904\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7737\
        );

    \I__903\ : Span4Mux_v
    port map (
            O => \N__7740\,
            I => \N__7734\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__7737\,
            I => \N__7731\
        );

    \I__901\ : Odrv4
    port map (
            O => \N__7734\,
            I => un5_visibley_ac0_11_0_1
        );

    \I__900\ : Odrv4
    port map (
            O => \N__7731\,
            I => un5_visibley_ac0_11_0_1
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__7726\,
            I => \N__7723\
        );

    \I__898\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7720\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__7720\,
            I => \un114_pixel_1_0_3__un1_beamylto9_3\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__7717\,
            I => \N__7714\
        );

    \I__895\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7711\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7705\
        );

    \I__893\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7702\
        );

    \I__892\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7697\
        );

    \I__891\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7697\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__7705\,
            I => \beamY_fastZ0Z_2\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__7702\,
            I => \beamY_fastZ0Z_2\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__7697\,
            I => \beamY_fastZ0Z_2\
        );

    \I__887\ : InMux
    port map (
            O => \N__7690\,
            I => \N__7684\
        );

    \I__886\ : InMux
    port map (
            O => \N__7689\,
            I => \N__7684\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__7684\,
            I => \N__7678\
        );

    \I__884\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7673\
        );

    \I__883\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7673\
        );

    \I__882\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7670\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__7678\,
            I => \N__7665\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__7673\,
            I => \N__7665\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__7670\,
            I => \N__7659\
        );

    \I__878\ : Span4Mux_h
    port map (
            O => \N__7665\,
            I => \N__7656\
        );

    \I__877\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7651\
        );

    \I__876\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7651\
        );

    \I__875\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7648\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__7659\,
            I => \beamYZ0Z_5\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__7656\,
            I => \beamYZ0Z_5\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__7651\,
            I => \beamYZ0Z_5\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__7648\,
            I => \beamYZ0Z_5\
        );

    \I__870\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7635\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__7638\,
            I => \N__7630\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__7635\,
            I => \N__7627\
        );

    \I__867\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7624\
        );

    \I__866\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7619\
        );

    \I__865\ : InMux
    port map (
            O => \N__7630\,
            I => \N__7619\
        );

    \I__864\ : Odrv12
    port map (
            O => \N__7627\,
            I => \beamY_fastZ0Z_3\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__7624\,
            I => \beamY_fastZ0Z_3\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__7619\,
            I => \beamY_fastZ0Z_3\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__7612\,
            I => \beamY_fast_RNIM4P7Z0Z_2_cascade_\
        );

    \I__860\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7601\
        );

    \I__859\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7601\
        );

    \I__858\ : InMux
    port map (
            O => \N__7607\,
            I => \N__7597\
        );

    \I__857\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7594\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7591\
        );

    \I__855\ : InMux
    port map (
            O => \N__7600\,
            I => \N__7585\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7580\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__7594\,
            I => \N__7580\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__7591\,
            I => \N__7577\
        );

    \I__851\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7574\
        );

    \I__850\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7569\
        );

    \I__849\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7569\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__7585\,
            I => \beamYZ0Z_6\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__7580\,
            I => \beamYZ0Z_6\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__7577\,
            I => \beamYZ0Z_6\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__7574\,
            I => \beamYZ0Z_6\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__7569\,
            I => \beamYZ0Z_6\
        );

    \I__843\ : InMux
    port map (
            O => \N__7558\,
            I => \N__7555\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__7555\,
            I => chessboardpixel_un174_pixel_0_1
        );

    \I__841\ : InMux
    port map (
            O => \N__7552\,
            I => \N__7549\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__7549\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0
        );

    \I__839\ : InMux
    port map (
            O => \N__7546\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__838\ : InMux
    port map (
            O => \N__7543\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5
        );

    \I__837\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7534\
        );

    \I__836\ : InMux
    port map (
            O => \N__7539\,
            I => \N__7534\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__7534\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8
        );

    \I__834\ : InMux
    port map (
            O => \N__7531\,
            I => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__832\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7522\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__7522\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHFZ0\
        );

    \I__830\ : InMux
    port map (
            O => \N__7519\,
            I => \N__7516\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__7516\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJZ0Z5\
        );

    \I__828\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7509\
        );

    \I__827\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7506\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__7509\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__7506\,
            I => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0\
        );

    \I__824\ : InMux
    port map (
            O => \N__7501\,
            I => \N__7498\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__7498\,
            I => \un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1Z0Z_1\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__7495\,
            I => \chessboardpixel_un200_pixel_0_1_cascade_\
        );

    \I__821\ : InMux
    port map (
            O => \N__7492\,
            I => \N__7489\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__7489\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__7486\,
            I => \N__7480\
        );

    \I__818\ : InMux
    port map (
            O => \N__7485\,
            I => \N__7477\
        );

    \I__817\ : InMux
    port map (
            O => \N__7484\,
            I => \N__7472\
        );

    \I__816\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7472\
        );

    \I__815\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7469\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__7477\,
            I => \beamY_i_2\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__7472\,
            I => \beamY_i_2\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__7469\,
            I => \beamY_i_2\
        );

    \I__811\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7456\
        );

    \I__810\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7456\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__7456\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81BZ0\
        );

    \I__808\ : InMux
    port map (
            O => \N__7453\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__806\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7444\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__7444\,
            I => \N__7441\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__7441\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEGZ0Z5\
        );

    \I__803\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7432\
        );

    \I__802\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7432\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__7432\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODGZ0\
        );

    \I__800\ : InMux
    port map (
            O => \N__7429\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3
        );

    \I__799\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7423\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__7423\,
            I => \N__7420\
        );

    \I__797\ : Odrv4
    port map (
            O => \N__7420\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87VZ0Z68\
        );

    \I__796\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7414\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__7414\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4JZ0\
        );

    \I__794\ : InMux
    port map (
            O => \N__7411\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__792\ : InMux
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__7399\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05UZ0Z8\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__7396\,
            I => \N__7392\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__7395\,
            I => \N__7388\
        );

    \I__787\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7377\
        );

    \I__786\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7377\
        );

    \I__785\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7377\
        );

    \I__784\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7377\
        );

    \I__783\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7374\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__7377\,
            I => \N__7371\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__7374\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__7371\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0\
        );

    \I__779\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7363\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__7363\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7
        );

    \I__777\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7357\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__7357\,
            I => \N__7354\
        );

    \I__775\ : Odrv4
    port map (
            O => \N__7354\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7
        );

    \I__774\ : InMux
    port map (
            O => \N__7351\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6
        );

    \I__773\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7339\
        );

    \I__772\ : InMux
    port map (
            O => \N__7347\,
            I => \N__7339\
        );

    \I__771\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7339\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__7339\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGKZ0\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__768\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7326\
        );

    \I__767\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7326\
        );

    \I__766\ : InMux
    port map (
            O => \N__7331\,
            I => \N__7323\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__7326\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__7323\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1\
        );

    \I__763\ : InMux
    port map (
            O => \N__7318\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4
        );

    \I__762\ : InMux
    port map (
            O => \N__7315\,
            I => \N__7312\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__7312\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\
        );

    \I__760\ : InMux
    port map (
            O => \N__7309\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5
        );

    \I__759\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7303\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__7303\,
            I => \beamY_RNIFJ0L_0Z0Z_8\
        );

    \I__757\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7297\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__7297\,
            I => \beamY_RNI19IJ_0Z0Z_9\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__7294\,
            I => \N__7290\
        );

    \I__754\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7280\
        );

    \I__753\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7280\
        );

    \I__752\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7280\
        );

    \I__751\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7277\
        );

    \I__750\ : InMux
    port map (
            O => \N__7287\,
            I => \N__7274\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__7280\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__7277\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__7274\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9\
        );

    \I__746\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7264\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__7264\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__7261\,
            I => \beamY_i_2_cascade_\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__7258\,
            I => \un114_pixel_1_0_3__chessboardpixel_un200_pixellto4Z0Z_1_cascade_\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__7255\,
            I => \chessboardpixel_un200_pixellt10_cascade_\
        );

    \I__741\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__7249\,
            I => un5_visibley_c6_0_0_0
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__7246\,
            I => \beamY_fast_RNI35GAZ0Z_2_cascade_\
        );

    \I__738\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7239\
        );

    \I__737\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7236\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__7239\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__7236\,
            I => \un21_beamy_cry_2_c_RNICOZ0Z83\
        );

    \I__734\ : InMux
    port map (
            O => \N__7231\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2
        );

    \I__733\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7225\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__7225\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2LZ0\
        );

    \I__731\ : InMux
    port map (
            O => \N__7222\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2
        );

    \I__730\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7216\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__7216\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO\
        );

    \I__728\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7210\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__7210\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RCZ0\
        );

    \I__726\ : InMux
    port map (
            O => \N__7207\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3
        );

    \I__725\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7200\
        );

    \I__724\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7197\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7200\,
            I => \un21_beamy_cry_6_c_RNIK4DZ0Z3\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__7197\,
            I => \un21_beamy_cry_6_c_RNIK4DZ0Z3\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__7192\,
            I => \N__7188\
        );

    \I__720\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7183\
        );

    \I__719\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7183\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__7183\,
            I => \beamY_fastZ0Z_7\
        );

    \I__717\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7177\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__7177\,
            I => \beamY_fastZ0Z_5\
        );

    \I__715\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7170\
        );

    \I__714\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7167\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__7170\,
            I => \un21_beamy_cry_1_c_RNIALZ0Z73\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__7167\,
            I => \un21_beamy_cry_1_c_RNIALZ0Z73\
        );

    \I__711\ : InMux
    port map (
            O => \N__7162\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2
        );

    \I__710\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7156\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__7156\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CRZ0Z2\
        );

    \I__708\ : InMux
    port map (
            O => \N__7153\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__7150\,
            I => \N__7147\
        );

    \I__706\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__7144\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGIZ0Z3\
        );

    \I__704\ : InMux
    port map (
            O => \N__7141\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__702\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__7132\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJZ0Z6874\
        );

    \I__700\ : InMux
    port map (
            O => \N__7129\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5
        );

    \I__699\ : InMux
    port map (
            O => \N__7126\,
            I => \N__7123\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__7123\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7
        );

    \I__697\ : InMux
    port map (
            O => \N__7120\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__7117\,
            I => \N__7114\
        );

    \I__695\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7111\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__7111\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__7108\,
            I => \N__7103\
        );

    \I__692\ : InMux
    port map (
            O => \N__7107\,
            I => \N__7098\
        );

    \I__691\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7089\
        );

    \I__690\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7089\
        );

    \I__689\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7089\
        );

    \I__688\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7089\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__7098\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__7089\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25\
        );

    \I__685\ : InMux
    port map (
            O => \N__7084\,
            I => \N__7081\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__7081\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7
        );

    \I__683\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7074\
        );

    \I__682\ : InMux
    port map (
            O => \N__7077\,
            I => \N__7071\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7074\,
            I => \N__7066\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__7071\,
            I => \N__7066\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__7066\,
            I => \un21_beamy_cry_4_c_RNIGUAZ0Z3\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__677\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__7057\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0
        );

    \I__675\ : InMux
    port map (
            O => \N__7054\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__673\ : InMux
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__7045\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICMZ0Z321\
        );

    \I__671\ : InMux
    port map (
            O => \N__7042\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3
        );

    \I__670\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7036\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__7036\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPMZ0Z1\
        );

    \I__668\ : InMux
    port map (
            O => \N__7033\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__7030\,
            I => \N__7027\
        );

    \I__666\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7024\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__7024\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KHZ0Z2\
        );

    \I__664\ : InMux
    port map (
            O => \N__7021\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5
        );

    \I__663\ : InMux
    port map (
            O => \N__7018\,
            I => \N__7015\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__7015\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7
        );

    \I__661\ : InMux
    port map (
            O => \N__7012\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__7009\,
            I => \N__7004\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__7008\,
            I => \N__7000\
        );

    \I__658\ : InMux
    port map (
            O => \N__7007\,
            I => \N__6996\
        );

    \I__657\ : InMux
    port map (
            O => \N__7004\,
            I => \N__6987\
        );

    \I__656\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6987\
        );

    \I__655\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6987\
        );

    \I__654\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6987\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__6996\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__6987\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92\
        );

    \I__651\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__6979\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_7
        );

    \I__649\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6973\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__6973\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0
        );

    \I__647\ : InMux
    port map (
            O => \N__6970\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6
        );

    \I__646\ : CascadeMux
    port map (
            O => \N__6967\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01_cascade_\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__6964\,
            I => \N__6961\
        );

    \I__644\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6958\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__6958\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0
        );

    \I__642\ : InMux
    port map (
            O => \N__6955\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2
        );

    \I__641\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6949\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__6949\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOLZ0\
        );

    \I__639\ : InMux
    port map (
            O => \N__6946\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__6943\,
            I => \N__6939\
        );

    \I__637\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6930\
        );

    \I__636\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6930\
        );

    \I__635\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6930\
        );

    \I__634\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6927\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__6930\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__6927\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__630\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6916\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__6916\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IGZ0Z1\
        );

    \I__628\ : InMux
    port map (
            O => \N__6913\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4
        );

    \I__627\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6907\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__6907\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__6904\,
            I => \N__6901\
        );

    \I__624\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6898\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__6898\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMGZ0Z1\
        );

    \I__622\ : InMux
    port map (
            O => \N__6895\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5
        );

    \I__621\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6889\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__6889\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7
        );

    \I__619\ : InMux
    port map (
            O => \N__6886\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6
        );

    \I__618\ : InMux
    port map (
            O => \N__6883\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6
        );

    \I__617\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6877\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__6877\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOGZ0Z53\
        );

    \I__615\ : InMux
    port map (
            O => \N__6874\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2
        );

    \I__614\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6868\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__6868\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOSZ0\
        );

    \I__612\ : InMux
    port map (
            O => \N__6865\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__6862\,
            I => \N__6859\
        );

    \I__610\ : InMux
    port map (
            O => \N__6859\,
            I => \N__6856\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__6856\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRSZ0\
        );

    \I__608\ : InMux
    port map (
            O => \N__6853\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__6850\,
            I => \N__6847\
        );

    \I__606\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6844\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__6844\,
            I => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LKZ0\
        );

    \I__604\ : InMux
    port map (
            O => \N__6841\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5
        );

    \I__603\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6835\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__6835\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_axb_7
        );

    \I__601\ : InMux
    port map (
            O => \N__6832\,
            I => un21_beamy_cry_5
        );

    \I__600\ : InMux
    port map (
            O => \N__6829\,
            I => un21_beamy_cry_6
        );

    \I__599\ : InMux
    port map (
            O => \N__6826\,
            I => un21_beamy_cry_7
        );

    \I__598\ : InMux
    port map (
            O => \N__6823\,
            I => \bfn_1_7_0_\
        );

    \I__597\ : InMux
    port map (
            O => \N__6820\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2
        );

    \I__596\ : InMux
    port map (
            O => \N__6817\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3
        );

    \I__595\ : InMux
    port map (
            O => \N__6814\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4
        );

    \I__594\ : InMux
    port map (
            O => \N__6811\,
            I => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5
        );

    \I__593\ : InMux
    port map (
            O => \N__6808\,
            I => un21_beamy_cry_1
        );

    \I__592\ : InMux
    port map (
            O => \N__6805\,
            I => un21_beamy_cry_2
        );

    \I__591\ : InMux
    port map (
            O => \N__6802\,
            I => un21_beamy_cry_3
        );

    \I__590\ : InMux
    port map (
            O => \N__6799\,
            I => un21_beamy_cry_4
        );

    \I__589\ : IoInMux
    port map (
            O => \N__6796\,
            I => \N__6793\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__6793\,
            I => \N__6790\
        );

    \I__587\ : Span4Mux_s1_h
    port map (
            O => \N__6790\,
            I => \N__6787\
        );

    \I__586\ : Span4Mux_h
    port map (
            O => \N__6787\,
            I => \N__6784\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__6784\,
            I => \N__6781\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__6781\,
            I => \Clock50MHz.PixelClock\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un8_beamx_cry_8,
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_6_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_10_0_\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un5_visiblex_cry_7,
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => un21_beamy_cry_8,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_7_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_8_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_4_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_11_0_\
        );

    \IN_MUX_bfv_9_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_8_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_10_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_10_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_7_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_9_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6796\,
            GLOBALBUFFEROUTPUT => \PixelClock_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \beamY_5_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7077\,
            lcout => \beamYZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11877\,
            ce => \N__11058\,
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un5_beamx_4_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7590\,
            in2 => \_gnd_net_\,
            in3 => \N__7663\,
            lcout => un1_beamy_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI6125_5_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101010101"
        )
    port map (
            in0 => \N__7664\,
            in1 => \N__12177\,
            in2 => \N__10632\,
            in3 => \N__8607\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBFP3_4_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__10595\,
            in1 => \N__12178\,
            in2 => \_gnd_net_\,
            in3 => \N__8608\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14760\,
            in2 => \N__15008\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => un21_beamy_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_1_c_RNIAL73_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12208\,
            in2 => \_gnd_net_\,
            in3 => \N__6808\,
            lcout => \un21_beamy_cry_1_c_RNIALZ0Z73\,
            ltout => OPEN,
            carryin => un21_beamy_cry_1,
            carryout => un21_beamy_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_2_c_RNICO83_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10631\,
            in2 => \_gnd_net_\,
            in3 => \N__6805\,
            lcout => \un21_beamy_cry_2_c_RNICOZ0Z83\,
            ltout => OPEN,
            carryin => un21_beamy_cry_2,
            carryout => un21_beamy_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_4_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10978\,
            in1 => \N__8620\,
            in2 => \_gnd_net_\,
            in3 => \N__6802\,
            lcout => \beamYZ0Z_4\,
            ltout => OPEN,
            carryin => un21_beamy_cry_3,
            carryout => un21_beamy_cry_4,
            clk => \N__11873\,
            ce => \N__11065\,
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_4_c_RNIGUA3_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7681\,
            in2 => \_gnd_net_\,
            in3 => \N__6799\,
            lcout => \un21_beamy_cry_4_c_RNIGUAZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_4,
            carryout => un21_beamy_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_6_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7600\,
            in2 => \_gnd_net_\,
            in3 => \N__6832\,
            lcout => \beamYZ0Z_6\,
            ltout => OPEN,
            carryin => un21_beamy_cry_5,
            carryout => un21_beamy_cry_6,
            clk => \N__11873\,
            ce => \N__11065\,
            sr => \_gnd_net_\
        );

    \un21_beamy_cry_6_c_RNIK4D3_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7809\,
            in2 => \_gnd_net_\,
            in3 => \N__6829\,
            lcout => \un21_beamy_cry_6_c_RNIK4DZ0Z3\,
            ltout => OPEN,
            carryin => un21_beamy_cry_6,
            carryout => un21_beamy_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_8_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7922\,
            in2 => \_gnd_net_\,
            in3 => \N__6826\,
            lcout => \beamYZ0Z_8\,
            ltout => OPEN,
            carryin => un21_beamy_cry_7,
            carryout => un21_beamy_cry_8,
            clk => \N__11873\,
            ce => \N__11065\,
            sr => \_gnd_net_\
        );

    \beamY_9_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10954\,
            in1 => \N__7852\,
            in2 => \_gnd_net_\,
            in3 => \N__6823\,
            lcout => \beamYZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11872\,
            ce => \N__11068\,
            sr => \_gnd_net_\
        );

    \beamY_7_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7203\,
            in2 => \_gnd_net_\,
            in3 => \N__10955\,
            lcout => \beamYZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11872\,
            ce => \N__11068\,
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12804\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOS_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7306\,
            in2 => \N__16402\,
            in3 => \N__6820\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNINGOSZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRS_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7228\,
            in2 => \N__16407\,
            in3 => \N__6817\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIKSRSZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LK_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7213\,
            in2 => \N__16403\,
            in3 => \N__6814\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI13LKZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI8C3M_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7288\,
            in1 => \N__6880\,
            in2 => \N__7336\,
            in3 => \N__6811\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6883\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_3_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12245\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOG53_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__7331\,
            in1 => \N__7332\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNIOGZ0Z53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_1_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9462\,
            in3 => \N__10891\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_c5_0_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOL_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7289\,
            in2 => \N__6964\,
            in3 => \N__6874\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNI5QOLZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IG1_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6871\,
            in2 => \N__7294\,
            in3 => \N__6865\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNI04IGZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMG1_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7293\,
            in2 => \N__6862\,
            in3 => \N__6853\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIUHMGZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNI70192_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6937\,
            in1 => \N__7267\,
            in2 => \N__6850\,
            in3 => \N__6841\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6970\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01\,
            ltout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5GZ0Z01_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIR5G01_0_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6967\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12805\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9535\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICM321_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6938\,
            in2 => \N__7063\,
            in3 => \N__6955\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNICMZ0Z321\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPM1_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6952\,
            in2 => \N__6943\,
            in3 => \N__6946\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIESPMZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KH2_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6942\,
            in2 => \N__6922\,
            in3 => \N__6913\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIA8KHZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI1RER4_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7007\,
            in1 => \N__6910\,
            in2 => \N__6904\,
            in3 => \N__6895\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6892\,
            in2 => \_gnd_net_\,
            in3 => \N__6886\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2LZ0Z92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9463\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHGR8_5_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__9537\,
            in1 => \N__9698\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => g0_2_0,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CR2_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6976\,
            in2 => \N__7008\,
            in3 => \N__7054\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_RNI57CRZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGI3_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7003\,
            in2 => \N__7051\,
            in3 => \N__7042\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGUGIZ0Z3\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJ6874_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7039\,
            in2 => \N__7009\,
            in3 => \N__7033\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIJZ0Z6874\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNI0RD4A_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7107\,
            in1 => \N__6982\,
            in2 => \N__7030\,
            in3 => \N__7021\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7018\,
            in2 => \_gnd_net_\,
            in3 => \N__7012\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6AZ0Z25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIO2L92_0_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6999\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9536\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un54_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8522\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEG5_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7102\,
            in2 => \N__7117\,
            in3 => \N__7162\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNI2AEGZ0Z5\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87V68_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7159\,
            in2 => \N__7108\,
            in3 => \N__7153\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNI87VZ0Z68\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05U8_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7106\,
            in2 => \N__7150\,
            in3 => \N__7141\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIK05UZ0Z8\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIE5N0K_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__7386\,
            in1 => \N__7084\,
            in2 => \N__7138\,
            in3 => \N__7129\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_axb_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDA_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7126\,
            in2 => \_gnd_net_\,
            in3 => \N__7120\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIMQPDAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9699\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIG6A25_0_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7101\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un61_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_5_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7078\,
            lcout => \beamY_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11880\,
            ce => \N__11057\,
            sr => \_gnd_net_\
        );

    \beamY_2_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7174\,
            lcout => \beamYZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11878\,
            ce => \N__11067\,
            sr => \_gnd_net_\
        );

    \beamY_3_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10974\,
            in2 => \_gnd_net_\,
            in3 => \N__7243\,
            lcout => \beamYZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11878\,
            ce => \N__11067\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIVDP7_7_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7911\,
            in1 => \N__7588\,
            in2 => \N__7192\,
            in3 => \N__7662\,
            lcout => un5_visibley_ac0_11_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_7_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__10975\,
            in1 => \N__7204\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11878\,
            ce => \N__11067\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIEP79_5_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7191\,
            in1 => \N__7180\,
            in2 => \_gnd_net_\,
            in3 => \N__7589\,
            lcout => un5_visibley_c6_0_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIP81D_7_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111110000"
        )
    port map (
            in0 => \N__8601\,
            in1 => \N__7994\,
            in2 => \N__7810\,
            in3 => \N__7955\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7173\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11875\,
            ce => \N__11066\,
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI35GA_0_2_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7708\,
            in1 => \N__7906\,
            in2 => \N__7638\,
            in3 => \N__8599\,
            lcout => un5_visibley_ac0_11_d,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNI35GA_2_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011100001111"
        )
    port map (
            in0 => \N__8600\,
            in1 => \N__7633\,
            in2 => \N__7923\,
            in3 => \N__7709\,
            lcout => OPEN,
            ltout => \beamY_fast_RNI35GAZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFJ0L_8_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__7252\,
            in1 => \_gnd_net_\,
            in2 => \N__7246\,
            in3 => \N__7910\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_3_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7242\,
            in2 => \_gnd_net_\,
            in3 => \N__10976\,
            lcout => \beamY_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11875\,
            ce => \N__11066\,
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_c_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12538\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_LUT4_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7231\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un26_sum_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI19IJ_9_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__7844\,
            in1 => \N__7758\,
            in2 => \_gnd_net_\,
            in3 => \N__7743\,
            lcout => chary_if_generate_plus_mult1_un33_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un8_beamylto4_0_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7634\,
            lcout => un5_visibley_c2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12654\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2L_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7300\,
            in2 => \N__16383\,
            in3 => \N__7222\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNIBT2LZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RC_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7219\,
            in2 => \N__16384\,
            in3 => \N__7207\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNIN1RCZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOI1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16355\,
            in2 => \_gnd_net_\,
            in3 => \N__7318\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4_c_RNICOIZ0Z1\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7315\,
            in2 => \_gnd_net_\,
            in3 => \N__7309\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVFZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFJ0L_0_8_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12655\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \beamY_RNIFJ0L_0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI19IJ_0_9_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12539\,
            lcout => \beamY_RNI19IJ_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un33_sum_cry_5_c_RNIPVF9_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7287\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un40_sum_i_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__7484\,
            in1 => \N__16401\,
            in2 => \_gnd_net_\,
            in3 => \N__12246\,
            lcout => \beamY_i_2\,
            ltout => \beamY_i_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_1_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010001000"
        )
    port map (
            in0 => \N__7461\,
            in1 => \N__7437\,
            in2 => \N__7261\,
            in3 => \N__7346\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__chessboardpixel_un200_pixellto4Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__chessboardpixel_un200_pixellto4_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001000000"
        )
    port map (
            in0 => \N__7347\,
            in1 => \N__15013\,
            in2 => \N__7258\,
            in3 => \N__7485\,
            lcout => OPEN,
            ltout => \chessboardpixel_un200_pixellt10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__chessboardpixel_un200_pixellto10_1_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000101"
        )
    port map (
            in0 => \N__7417\,
            in1 => \N__7492\,
            in2 => \N__7255\,
            in3 => \N__7348\,
            lcout => OPEN,
            ltout => \chessboardpixel_un200_pixel_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__Pixel_3_sqmuxa_0_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12118\,
            in2 => \N__7495\,
            in3 => \N__7558\,
            lcout => \un114_pixel_1_0_3__Pixel_3_sqmuxaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIMR0FR_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__7462\,
            in1 => \N__7483\,
            in2 => \_gnd_net_\,
            in3 => \N__7438\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un1_rem_adjust_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7486\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81B_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7552\,
            in2 => \N__7395\,
            in3 => \N__7453\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_RNIDK81BZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODG_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7391\,
            in2 => \N__7450\,
            in3 => \N__7429\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI97ODGZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4J_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7426\,
            in2 => \N__7396\,
            in3 => \N__7411\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIG6A4JZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7366\,
            in2 => \N__7408\,
            in3 => \N__7387\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_7,
            ltout => OPEN,
            carryin => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGK_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7360\,
            in2 => \_gnd_net_\,
            in3 => \N__7351\,
            lcout => \chessboardpixel_un178_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNI2EAGKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001010010010"
        )
    port map (
            in0 => \N__7501\,
            in1 => \N__7513\,
            in2 => \N__7528\,
            in3 => \N__11544\,
            lcout => chessboardpixel_un174_pixel_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8523\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un68_sum_i_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11547\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJ5_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7539\,
            in2 => \N__9043\,
            in3 => \N__7546\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI3JJZ0Z5\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAEC_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8203\,
            in2 => \N__8248\,
            in3 => \N__7543\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5_c_RNIDLAECZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8202\,
            in1 => \N__7540\,
            in2 => \N__8233\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHF_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8218\,
            in2 => \_gnd_net_\,
            in3 => \N__7531\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNIL0DHFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1_1_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100010101"
        )
    port map (
            in0 => \N__7519\,
            in1 => \N__7512\,
            in2 => \N__13612\,
            in3 => \N__11548\,
            lcout => \un114_pixel_1_0_3__chessboardpixel_un174_pixellto10_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKHPCA1_4_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9765\,
            in1 => \N__9298\,
            in2 => \_gnd_net_\,
            in3 => \N__9933\,
            lcout => \beamY_RNIKHPCA1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNISKOB_5_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010010101"
        )
    port map (
            in0 => \N__7608\,
            in1 => \N__8641\,
            in2 => \N__8008\,
            in3 => \N__7682\,
            lcout => chessboardpixel_un178_pixel_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un1_beamylto9_0_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10641\,
            in2 => \_gnd_net_\,
            in3 => \N__7825\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un1_beamylto9Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un1_beamylto9_3_0_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110000"
        )
    port map (
            in0 => \N__14994\,
            in1 => \N__12216\,
            in2 => \N__7768\,
            in3 => \N__8642\,
            lcout => \un114_pixel_1_0_3__un1_beamylto9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_1_3_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10640\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12215\,
            lcout => un4_beamylt6,
            ltout => \un4_beamylt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_beamylto6_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__7683\,
            in1 => \N__7609\,
            in2 => \N__7765\,
            in3 => \N__8643\,
            lcout => un4_beamylt8_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIDO3I_9_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110101010101"
        )
    port map (
            in0 => \N__7871\,
            in1 => \N__7823\,
            in2 => \N__8038\,
            in3 => \N__7924\,
            lcout => \beamY_RNIDO3IZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGSI81_9_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001100000"
        )
    port map (
            in0 => \N__7870\,
            in1 => \N__7762\,
            in2 => \N__12685\,
            in3 => \N__7747\,
            lcout => chary_if_generate_plus_mult1_un40_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un1_beamylto9_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7872\,
            in1 => \N__7978\,
            in2 => \N__7726\,
            in3 => \N__7925\,
            lcout => un1_beamylto9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIM4P7_2_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__8629\,
            in1 => \N__7606\,
            in2 => \N__7717\,
            in3 => \N__7689\,
            lcout => OPEN,
            ltout => \beamY_fast_RNIM4P7Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_fast_RNIJP9E_3_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__7690\,
            in1 => \N__7639\,
            in2 => \N__7612\,
            in3 => \N__7607\,
            lcout => un5_visibley_c5,
            ltout => \un5_visibley_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI0A5O1_7_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110111"
        )
    port map (
            in0 => \N__7824\,
            in1 => \N__12665\,
            in2 => \N__8029\,
            in3 => \N__12581\,
            lcout => chary_if_generate_plus_mult1_un40_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un5_beamx_5_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7819\,
            in1 => \N__15007\,
            in2 => \N__8659\,
            in3 => \N__7874\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un5_beamxZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un5_beamx_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8645\,
            in1 => \N__7977\,
            in2 => \N__8026\,
            in3 => \N__7939\,
            lcout => un5_beamx_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_1_0_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7875\,
            in2 => \_gnd_net_\,
            in3 => \N__7938\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__g0_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7976\,
            in1 => \N__8563\,
            in2 => \N__8023\,
            in3 => \N__7818\,
            lcout => un1_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_beamylto9_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__7816\,
            in1 => \N__7873\,
            in2 => \N__8020\,
            in3 => \N__7936\,
            lcout => un4_beamy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un8_beamylto9_1_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__8004\,
            in1 => \N__7975\,
            in2 => \_gnd_net_\,
            in3 => \N__8644\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un8_beamylto9Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un8_beamylto9_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7937\,
            in1 => \N__7876\,
            in2 => \N__7828\,
            in3 => \N__7817\,
            lcout => un8_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc3_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9764\,
            in1 => \N__8064\,
            in2 => \N__8548\,
            in3 => \N__8157\,
            lcout => if_generate_plus_mult1_un75_sum_axbxc3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un54_sum_c5_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001001100100"
        )
    port map (
            in0 => \N__12816\,
            in1 => \N__12687\,
            in2 => \N__9460\,
            in3 => \N__12591\,
            lcout => \row_1_if_generate_plus_mult1_un54_sum_cZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axbxc5_1_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000110000111"
        )
    port map (
            in0 => \N__8080\,
            in1 => \N__8050\,
            in2 => \N__12417\,
            in3 => \N__12437\,
            lcout => \row_1_if_generate_plus_mult1_un82_sum_axbxc5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_c5_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101110000010"
        )
    port map (
            in0 => \N__8079\,
            in1 => \N__8065\,
            in2 => \N__8158\,
            in3 => \N__8049\,
            lcout => \row_1_if_generate_plus_mult1_un75_sum_cZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_c4_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000011110110"
        )
    port map (
            in0 => \N__8063\,
            in1 => \N__8153\,
            in2 => \N__8547\,
            in3 => \N__9763\,
            lcout => \row_1_if_generate_plus_mult1_un75_sum_cZ0Z4\,
            ltout => \row_1_if_generate_plus_mult1_un75_sum_cZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101001"
        )
    port map (
            in0 => \N__12410\,
            in1 => \N__8048\,
            in2 => \N__8071\,
            in3 => \N__12436\,
            lcout => if_generate_plus_mult1_un75_sum_axbxc5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_c4_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__8131\,
            in1 => \N__10877\,
            in2 => \_gnd_net_\,
            in3 => \N__9445\,
            lcout => OPEN,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_cZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_1_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10878\,
            in1 => \N__8125\,
            in2 => \N__8068\,
            in3 => \N__12721\,
            lcout => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1\,
            ltout => \row_1_if_generate_plus_mult1_un68_sum_axbxc5Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc5_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8053\,
            in3 => \N__8152\,
            lcout => if_generate_plus_mult1_un68_sum_axbxc5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_axbxc3_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__9762\,
            in1 => \N__12722\,
            in2 => \_gnd_net_\,
            in3 => \N__9591\,
            lcout => if_generate_plus_mult1_un68_sum_axbxc3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un54_sum_axbxc3_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100111010010"
        )
    port map (
            in0 => \N__12812\,
            in1 => \N__12679\,
            in2 => \N__9461\,
            in3 => \N__12592\,
            lcout => if_generate_plus_mult1_un54_sum_axbxc3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_c5_0_ns_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111001011000"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__8095\,
            in2 => \N__8170\,
            in3 => \N__9761\,
            lcout => row_1_if_generate_plus_mult1_un68_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9449\,
            in1 => \N__10883\,
            in2 => \_gnd_net_\,
            in3 => \N__9571\,
            lcout => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_axbxc5_1_0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100111011011"
        )
    port map (
            in0 => \N__12811\,
            in1 => \N__12689\,
            in2 => \N__12599\,
            in3 => \N__9448\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0\,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_axbxc5_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_axbxc5_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8110\,
            in2 => \N__8134\,
            in3 => \N__10882\,
            lcout => if_generate_plus_mult1_un61_sum_axbxc5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_5_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10879\,
            in1 => \N__9570\,
            in2 => \_gnd_net_\,
            in3 => \N__9446\,
            lcout => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5\,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_ac0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_7_0_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101010"
        )
    port map (
            in0 => \N__8089\,
            in1 => \N__8124\,
            in2 => \N__8113\,
            in3 => \N__10880\,
            lcout => row_1_if_generate_plus_mult1_un61_sum_c5,
            ltout => \row_1_if_generate_plus_mult1_un61_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un68_sum_c5_0_bm_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010100101"
        )
    port map (
            in0 => \N__10881\,
            in1 => \_gnd_net_\,
            in2 => \N__8104\,
            in3 => \N__8101\,
            lcout => if_generate_plus_mult1_un68_sum_c5_0_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un61_sum_ac0_7_c_0_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010010010"
        )
    port map (
            in0 => \N__12810\,
            in1 => \N__12688\,
            in2 => \N__12598\,
            in3 => \N__9447\,
            lcout => row_1_if_generate_plus_mult1_un61_sum_ac0_7_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11656\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_11_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KC4_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8184\,
            in2 => \N__9052\,
            in3 => \N__8236\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIN6KCZ0Z4\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGS6_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13957\,
            in2 => \N__13915\,
            in3 => \N__8221\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI6HGSZ0Z6\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI88ODF_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8201\,
            in1 => \N__8185\,
            in2 => \N__13945\,
            in3 => \N__8209\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un75_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3U7_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13930\,
            in2 => \_gnd_net_\,
            in3 => \N__8206\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIBQ3UZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13911\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_cry_1_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8263\,
            in2 => \N__8350\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => counter_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNO_0_2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8320\,
            in2 => \_gnd_net_\,
            in3 => \N__8176\,
            lcout => counter_30,
            ltout => OPEN,
            carryin => counter_cry_1,
            carryout => counter_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNO_0_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8366\,
            in2 => \_gnd_net_\,
            in3 => \N__8173\,
            lcout => counter_29,
            ltout => OPEN,
            carryin => counter_cry_2,
            carryout => counter_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNO_0_4_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8937\,
            in2 => \_gnd_net_\,
            in3 => \N__8293\,
            lcout => counter_28,
            ltout => OPEN,
            carryin => counter_cry_3,
            carryout => counter_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNO_0_5_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9021\,
            in2 => \_gnd_net_\,
            in3 => \N__8290\,
            lcout => counter_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNI6R5D_0_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8264\,
            in1 => \N__8368\,
            in2 => \N__8349\,
            in3 => \N__8319\,
            lcout => slaveselect_1_0_4,
            ltout => \slaveselect_1_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIVUOJ_5_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__8938\,
            in1 => \_gnd_net_\,
            in2 => \N__8287\,
            in3 => \N__9022\,
            lcout => un3_slaveselect,
            ltout => \un3_slaveselect_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_2_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011000100"
        )
    port map (
            in0 => \N__8900\,
            in1 => \N__8284\,
            in2 => \N__8278\,
            in3 => \N__8858\,
            lcout => \counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_3_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010100000000"
        )
    port map (
            in0 => \N__8851\,
            in1 => \N__8971\,
            in2 => \N__8911\,
            in3 => \N__8275\,
            lcout => \counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNO_0_1_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__8348\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8265\,
            lcout => OPEN,
            ltout => \counter_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_1_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010110000"
        )
    port map (
            in0 => \N__8970\,
            in1 => \N__8907\,
            in2 => \N__8269\,
            in3 => \N__8852\,
            lcout => \counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_0_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000101"
        )
    port map (
            in0 => \N__8850\,
            in1 => \N__8969\,
            in2 => \N__8910\,
            in3 => \N__8266\,
            lcout => \counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIKUI6_1_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8367\,
            in2 => \_gnd_net_\,
            in3 => \N__8347\,
            lcout => OPEN,
            ltout => \un1_counterlto3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNINHFG_2_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__8939\,
            in1 => \N__9023\,
            in2 => \N__8323\,
            in3 => \N__8318\,
            lcout => un1_counter_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIS857F2_4_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9934\,
            in1 => \N__10045\,
            in2 => \N__9783\,
            in3 => \N__9296\,
            lcout => OPEN,
            ltout => \g0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJU3OQ8_4_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001101001"
        )
    port map (
            in0 => \N__9361\,
            in1 => \N__9859\,
            in2 => \N__8302\,
            in3 => \N__9257\,
            lcout => g0_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUAPPF4_0_3_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110110001110"
        )
    port map (
            in0 => \N__10048\,
            in1 => \N__8546\,
            in2 => \N__9782\,
            in3 => \N__8299\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_1_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010000001"
        )
    port map (
            in0 => \N__8434\,
            in1 => \N__9081\,
            in2 => \N__8377\,
            in3 => \N__9358\,
            lcout => chary_if_generate_plus_mult1_un68_sum_0_0_0_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2TEJF4_0_4_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__10046\,
            in1 => \N__9846\,
            in2 => \_gnd_net_\,
            in3 => \N__9256\,
            lcout => chary_if_generate_plus_mult1_un61_sum_0_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHUG2_0_3_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10662\,
            in2 => \_gnd_net_\,
            in3 => \N__12247\,
            lcout => un5_visibley_0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIQ53PA3_4_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9845\,
            in2 => \_gnd_net_\,
            in3 => \N__9255\,
            lcout => chary_if_generate_plus_mult1_un61_sum_c5,
            ltout => \chary_if_generate_plus_mult1_un61_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIUAPPF4_3_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101110110010"
        )
    port map (
            in0 => \N__8443\,
            in1 => \N__9770\,
            in2 => \N__8437\,
            in3 => \N__10047\,
            lcout => chary_if_generate_plus_mult1_un68_sum_c4_0,
            ltout => \chary_if_generate_plus_mult1_un68_sum_c4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKP1Q9A_5_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001001110001"
        )
    port map (
            in0 => \N__8401\,
            in1 => \N__8433\,
            in2 => \N__8425\,
            in3 => \N__9923\,
            lcout => OPEN,
            ltout => \g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIBLQCVR_2_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001101001"
        )
    port map (
            in0 => \N__8422\,
            in1 => \N__9322\,
            in2 => \N__8416\,
            in3 => \N__12248\,
            lcout => g2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIV142B4_3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101101001"
        )
    port map (
            in0 => \N__9910\,
            in1 => \N__9348\,
            in2 => \N__9297\,
            in3 => \N__10642\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un75_sum_c5_N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICECPQ8_4_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011100010"
        )
    port map (
            in0 => \N__8413\,
            in1 => \N__9190\,
            in2 => \N__8404\,
            in3 => \N__8647\,
            lcout => chary_if_generate_plus_mult1_un75_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFJKLC_0_5_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9720\,
            in1 => \N__10085\,
            in2 => \N__9638\,
            in3 => \N__9545\,
            lcout => g0_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKHPCA1_5_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10086\,
            in1 => \N__9630\,
            in2 => \N__8395\,
            in3 => \N__9911\,
            lcout => chary_if_generate_plus_mult1_un61_sum_1_0_1_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI44RHC_5_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9626\,
            in1 => \N__10084\,
            in2 => \_gnd_net_\,
            in3 => \N__9542\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNINITP61_5_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011010100"
        )
    port map (
            in0 => \N__9544\,
            in1 => \N__10135\,
            in2 => \N__9739\,
            in3 => \N__9909\,
            lcout => OPEN,
            ltout => \beamY_RNINITP61Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITFRN03_5_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9137\,
            in2 => \N__8488\,
            in3 => \N__8485\,
            lcout => \beamY_RNITFRN03Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNINITP61_1_5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100101011"
        )
    port map (
            in0 => \N__9543\,
            in1 => \N__10134\,
            in2 => \N__9738\,
            in3 => \N__9908\,
            lcout => \beamY_RNINITP61_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIIIGJ2_0_9_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101001011110"
        )
    port map (
            in0 => \N__8478\,
            in1 => \N__9403\,
            in2 => \N__12809\,
            in3 => \N__9803\,
            lcout => chary_if_generate_plus_mult1_un47_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIIIGJ2_9_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110000111001"
        )
    port map (
            in0 => \N__12792\,
            in1 => \N__8479\,
            in2 => \N__9816\,
            in3 => \N__9427\,
            lcout => chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0,
            ltout => \chary_if_generate_plus_mult1_un54_sum_axbxc5_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI14TP8_7_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8701\,
            in1 => \N__8467\,
            in2 => \N__8470\,
            in3 => \N__8458\,
            lcout => chary_if_generate_plus_mult1_un54_sum_axbxc5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITKMQ1_9_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011001"
        )
    port map (
            in0 => \N__9808\,
            in1 => \N__12670\,
            in2 => \_gnd_net_\,
            in3 => \N__12584\,
            lcout => chary_if_generate_plus_mult1_un47_sum_axbxc5_2,
            ltout => \chary_if_generate_plus_mult1_un47_sum_axbxc5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIB65I6_7_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8700\,
            in1 => \N__8457\,
            in2 => \N__8461\,
            in3 => \N__9404\,
            lcout => chary_if_generate_plus_mult1_un54_sum_axb3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITURI3_7_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110010110"
        )
    port map (
            in0 => \N__8455\,
            in1 => \N__12666\,
            in2 => \N__9815\,
            in3 => \N__12582\,
            lcout => \beamY_RNITURI3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNITURI3_0_7_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__12583\,
            in1 => \N__8456\,
            in2 => \N__12686\,
            in3 => \N__9804\,
            lcout => OPEN,
            ltout => \beamY_RNITURI3_0Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNICG8P9_7_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8699\,
            in2 => \N__8689\,
            in3 => \N__8686\,
            lcout => \beamY_RNICG8P9Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un15_beamy_2_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8554\,
            in1 => \N__8680\,
            in2 => \N__10237\,
            in3 => \N__8674\,
            lcout => \un114_pixel_1_0_3__un15_beamyZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un3_beamx_2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10746\,
            in2 => \_gnd_net_\,
            in3 => \N__10281\,
            lcout => un1_beamx_2,
            ltout => \un1_beamx_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un15_beamy_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001100"
        )
    port map (
            in0 => \N__8755\,
            in1 => \N__8668\,
            in2 => \N__8662\,
            in3 => \N__10322\,
            lcout => un15_beamy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un5_beamx_3_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__14634\,
            in1 => \N__10667\,
            in2 => \_gnd_net_\,
            in3 => \N__12253\,
            lcout => \un114_pixel_1_0_3__un5_beamxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_1_3_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__12254\,
            in1 => \N__10668\,
            in2 => \N__15016\,
            in3 => \N__8646\,
            lcout => \un114_pixel_1_0_3__g0_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un18_beamylto9_2_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10273\,
            in1 => \N__10312\,
            in2 => \N__10747\,
            in3 => \N__10364\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un18_beamylto9Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un18_beamylto9_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__10188\,
            in1 => \N__10397\,
            in2 => \N__8557\,
            in3 => \N__10448\,
            lcout => un18_beamylt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_1_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000110101"
        )
    port map (
            in0 => \N__12251\,
            in1 => \N__8545\,
            in2 => \N__8749\,
            in3 => \N__10663\,
            lcout => \row_1_if_generate_plus_mult1_un82_sum_ac0_7_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un13_beamylto6_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010011"
        )
    port map (
            in0 => \N__10449\,
            in1 => \N__10365\,
            in2 => \N__10411\,
            in3 => \N__10189\,
            lcout => un13_beamylt7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_axb4_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12438\,
            in1 => \N__8736\,
            in2 => \N__12465\,
            in3 => \N__12406\,
            lcout => OPEN,
            ltout => \row_1_if_generate_plus_mult1_un82_sum_axb4_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un82_sum_ac0_7_0_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000100"
        )
    port map (
            in0 => \N__8748\,
            in1 => \N__8737\,
            in2 => \N__8725\,
            in3 => \N__8722\,
            lcout => row_1_if_generate_plus_mult1_un82_sum_c5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un8_beamx_cry_1_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10550\,
            in2 => \N__12024\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => un8_beamx_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_2_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10518\,
            in2 => \_gnd_net_\,
            in3 => \N__8716\,
            lcout => \beamXZ0Z_2\,
            ltout => OPEN,
            carryin => un8_beamx_cry_1,
            carryout => un8_beamx_cry_2,
            clk => \N__11874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10486\,
            in2 => \_gnd_net_\,
            in3 => \N__8713\,
            lcout => \beamXZ0Z_3\,
            ltout => OPEN,
            carryin => un8_beamx_cry_2,
            carryout => un8_beamx_cry_3,
            clk => \N__11874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_4_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11040\,
            in1 => \N__10451\,
            in2 => \_gnd_net_\,
            in3 => \N__8710\,
            lcout => \beamXZ0Z_4\,
            ltout => OPEN,
            carryin => un8_beamx_cry_3,
            carryout => un8_beamx_cry_4,
            clk => \N__11874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_5_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10414\,
            in2 => \_gnd_net_\,
            in3 => \N__8707\,
            lcout => \beamXZ0Z_5\,
            ltout => OPEN,
            carryin => un8_beamx_cry_4,
            carryout => un8_beamx_cry_5,
            clk => \N__11874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_6_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10367\,
            in2 => \_gnd_net_\,
            in3 => \N__8704\,
            lcout => \beamXZ0Z_6\,
            ltout => OPEN,
            carryin => un8_beamx_cry_5,
            carryout => un8_beamx_cry_6,
            clk => \N__11874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_7_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10321\,
            in2 => \_gnd_net_\,
            in3 => \N__8779\,
            lcout => \beamXZ0Z_7\,
            ltout => OPEN,
            carryin => un8_beamx_cry_6,
            carryout => un8_beamx_cry_7,
            clk => \N__11874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_8_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10277\,
            in2 => \_gnd_net_\,
            in3 => \N__8776\,
            lcout => \beamXZ0Z_8\,
            ltout => OPEN,
            carryin => un8_beamx_cry_7,
            carryout => un8_beamx_cry_8,
            clk => \N__11874\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_9_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10742\,
            in2 => \_gnd_net_\,
            in3 => \N__8773\,
            lcout => \beamXZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => un8_beamx_cry_9,
            clk => \N__11879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_10_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__10231\,
            in1 => \N__11042\,
            in2 => \_gnd_net_\,
            in3 => \N__8770\,
            lcout => \beamXZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8V_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10174\,
            in2 => \_gnd_net_\,
            in3 => \N__10175\,
            lcout => \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNI2R8VZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_1_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10551\,
            in2 => \_gnd_net_\,
            in3 => \N__12002\,
            lcout => \beamXZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11879\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1_2_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110101001011"
        )
    port map (
            in0 => \N__12723\,
            in1 => \N__9784\,
            in2 => \N__8767\,
            in3 => \N__9592\,
            lcout => \row_1_if_generate_plus_mult1_un75_sum_axbxc5_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__N_204_0_i_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16155\,
            in3 => \N__12937\,
            lcout => \N_204_0_i\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => charx_if_generate_plus_mult1_un19_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_LUT4_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8758\,
            lcout => \charx_if_generate_plus_mult1_un19_sum_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_0_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13872\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_0_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11649\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nCS1_1_RNO_0_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__9024\,
            in1 => \N__8893\,
            in2 => \N__8940\,
            in3 => \N__9000\,
            lcout => \nCS1_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_5_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000001100"
        )
    port map (
            in0 => \N__8968\,
            in1 => \N__9031\,
            in2 => \N__8860\,
            in3 => \N__8898\,
            lcout => \counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \slaveselect_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8894\,
            in1 => \N__8854\,
            in2 => \_gnd_net_\,
            in3 => \N__8966\,
            lcout => \slaveselectZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_RNIQHKU_5_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__9025\,
            in1 => \N__8899\,
            in2 => \N__8941\,
            in3 => \N__9001\,
            lcout => un1_slaveselect_1_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \counter_4_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010100000000"
        )
    port map (
            in0 => \N__8853\,
            in1 => \N__8967\,
            in2 => \N__8909\,
            in3 => \N__8947\,
            lcout => \counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14327\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \nCS1_1_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__8802\,
            in1 => \N__8908\,
            in2 => \_gnd_net_\,
            in3 => \N__8859\,
            lcout => \nCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14328\,
            ce => 'H',
            sr => \N__8791\
        );

    \un114_pixel_1_0_3__g0_8_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000010010"
        )
    port map (
            in0 => \N__9360\,
            in1 => \N__9088\,
            in2 => \N__9112\,
            in3 => \N__12250\,
            lcout => font_un28_pixel_0_0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2TEJF4_4_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__10043\,
            in1 => \N__9857\,
            in2 => \_gnd_net_\,
            in3 => \N__9254\,
            lcout => \beamY_RNI2TEJF4Z0Z_4\,
            ltout => \beamY_RNI2TEJF4Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_8_1_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010000001"
        )
    port map (
            in0 => \N__9221\,
            in1 => \N__9163\,
            in2 => \N__9115\,
            in3 => \N__10664\,
            lcout => \un114_pixel_1_0_3__g0_8Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKHPCA1_0_4_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9769\,
            in1 => \N__9295\,
            in2 => \_gnd_net_\,
            in3 => \N__9932\,
            lcout => chary_if_generate_plus_mult1_un61_sum_0_3,
            ltout => \chary_if_generate_plus_mult1_un61_sum_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_10_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10044\,
            in2 => \N__9103\,
            in3 => \N__9359\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__g0_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_3_0_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011100001"
        )
    port map (
            in0 => \N__9259\,
            in1 => \N__9858\,
            in2 => \N__9100\,
            in3 => \N__9325\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__g0_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_9_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011111100001"
        )
    port map (
            in0 => \N__9097\,
            in1 => \N__9186\,
            in2 => \N__9091\,
            in3 => \N__9162\,
            lcout => chary_if_generate_plus_mult1_un75_sum_i_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_6_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110001101001"
        )
    port map (
            in0 => \N__9855\,
            in1 => \N__10035\,
            in2 => \N__9952\,
            in3 => \N__9258\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__g0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_5_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9082\,
            in2 => \N__9070\,
            in3 => \N__9323\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__g0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_0_1_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101101111110"
        )
    port map (
            in0 => \N__9067\,
            in1 => \N__9061\,
            in2 => \N__9055\,
            in3 => \N__10665\,
            lcout => \un114_pixel_1_0_3__N_5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIH9THAD_4_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111010000001"
        )
    port map (
            in0 => \N__9184\,
            in1 => \N__9159\,
            in2 => \N__9226\,
            in3 => \N__9357\,
            lcout => \beamY_RNIH9THADZ0Z_4\,
            ltout => \beamY_RNIH9THADZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIHHB5F01_4_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9324\,
            in1 => \N__9196\,
            in2 => \N__9301\,
            in3 => \N__9161\,
            lcout => \beamY_RNIHHB5F01Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI3SPGT1_4_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001000000"
        )
    port map (
            in0 => \N__9139\,
            in1 => \N__9282\,
            in2 => \N__9781\,
            in3 => \N__9906\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_7_d,
            ltout => \chary_if_generate_plus_mult1_un61_sum_ac0_7_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIME80Q5_4_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__9856\,
            in1 => \N__9222\,
            in2 => \N__9199\,
            in3 => \N__10034\,
            lcout => chary_if_generate_plus_mult1_un68_sum_axb4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKP1Q9A_0_5_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100010000001"
        )
    port map (
            in0 => \N__9185\,
            in1 => \N__9160\,
            in2 => \N__9604\,
            in3 => \N__9907\,
            lcout => g1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFA04J_5_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9539\,
            in1 => \N__9479\,
            in2 => \N__9639\,
            in3 => \N__10083\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGS0LB_5_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110100"
        )
    port map (
            in0 => \N__10082\,
            in1 => \N__9538\,
            in2 => \N__10111\,
            in3 => \N__9450\,
            lcout => \beamY_RNIGS0LBZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNINITP61_0_5_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100101011"
        )
    port map (
            in0 => \N__9541\,
            in1 => \N__10138\,
            in2 => \N__9760\,
            in3 => \N__9924\,
            lcout => OPEN,
            ltout => \g0_0_x2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVC6VP1_3_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9138\,
            in2 => \N__9118\,
            in3 => \N__10658\,
            lcout => g0_0_x2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIC02EA1_2_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__9721\,
            in1 => \N__9823\,
            in2 => \N__9931\,
            in3 => \N__12249\,
            lcout => g0_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIARUFB_5_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__10109\,
            in1 => \N__10081\,
            in2 => \_gnd_net_\,
            in3 => \N__9451\,
            lcout => OPEN,
            ltout => \beamY_RNIARUFBZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI5U4NT_5_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9478\,
            in2 => \N__9943\,
            in3 => \N__9940\,
            lcout => chary_if_generate_plus_mult1_un54_sum_c5,
            ltout => \chary_if_generate_plus_mult1_un54_sum_c5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIN998D1_5_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110101010"
        )
    port map (
            in0 => \N__9480\,
            in1 => \N__10136\,
            in2 => \N__9862\,
            in3 => \N__9540\,
            lcout => chary_if_generate_plus_mult1_un61_sum_ac0_7_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI44RHC_0_5_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__9588\,
            in1 => \N__9634\,
            in2 => \_gnd_net_\,
            in3 => \N__10089\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axb3_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2MTA1_9_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__9817\,
            in1 => \N__9458\,
            in2 => \_gnd_net_\,
            in3 => \N__12791\,
            lcout => \beamY_RNI2MTA1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIFJKLC_5_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__10090\,
            in1 => \N__9780\,
            in2 => \N__9640\,
            in3 => \N__9589\,
            lcout => g0_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPC8SG_5_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__10087\,
            in1 => \N__9587\,
            in2 => \N__9484\,
            in3 => \N__9459\,
            lcout => OPEN,
            ltout => \chary_if_generate_plus_mult1_un54_sum_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI8NBQ41_5_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100101101010"
        )
    port map (
            in0 => \N__10137\,
            in1 => \N__10110\,
            in2 => \N__10093\,
            in3 => \N__10088\,
            lcout => chary_if_generate_plus_mult1_un61_sum_axbxc5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un3_beamx_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__10198\,
            in1 => \N__9996\,
            in2 => \N__10329\,
            in3 => \N__10412\,
            lcout => un3_beamx_0,
            ltout => \un3_beamx_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_0_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10970\,
            in2 => \N__10000\,
            in3 => \N__14641\,
            lcout => \beamYZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJPPPPD1_3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__12291\,
            in1 => \N__10666\,
            in2 => \N__10690\,
            in3 => \N__12252\,
            lcout => chary_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HSyncZ0_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__10236\,
            in1 => \N__9997\,
            in2 => \N__10330\,
            in3 => \N__10243\,
            lcout => \HSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11881\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15093\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIG328_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10144\,
            in2 => \_gnd_net_\,
            in3 => \N__9973\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_1_c_RNIGZ0Z328\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HL_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16364\,
            in2 => \N__10153\,
            in3 => \N__9970\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_2_c_RNI16HLZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_3_c_RNIMVPQ1_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11229\,
            in1 => \N__10180\,
            in2 => \N__9967\,
            in3 => \N__9955\,
            lcout => charx_if_generate_plus_mult1_un33_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un26_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un26_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10246\,
            lcout => \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISUZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un1_beamxlto6_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10413\,
            in1 => \N__10452\,
            in2 => \N__10492\,
            in3 => \N__10368\,
            lcout => un1_beamxlt10_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un3_beamx_5_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10549\,
            in1 => \N__10517\,
            in2 => \N__10235\,
            in3 => \N__10450\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un3_beamxZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un3_beamx_7_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10485\,
            in1 => \N__10366\,
            in2 => \N__10201\,
            in3 => \N__11989\,
            lcout => \un114_pixel_1_0_3__un3_beamxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_4_0_15__un13_beamylto3_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__10516\,
            in1 => \N__10548\,
            in2 => \N__10491\,
            in3 => \N__11988\,
            lcout => un18_beamylt4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamX_0_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11041\,
            lcout => \beamXZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11876\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKF_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10179\,
            lcout => \charx_if_generate_plus_mult1_un19_sum_cry_1_c_RNIHDKFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_N_575_i_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11645\,
            lcout => \N_575_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16156\,
            lcout => charx_if_generate_plus_mult1_un19_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12003\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_10_0_\,
            carryout => un5_visiblex_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_0_c_RNIHKT1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10552\,
            in3 => \N__10522\,
            lcout => charx_if_generate_plus_mult1_un75_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_0,
            carryout => un5_visiblex_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10519\,
            in3 => \N__10495\,
            lcout => charx_if_generate_plus_mult1_un68_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_1,
            carryout => un5_visiblex_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16394\,
            in2 => \N__10490\,
            in3 => \N__10456\,
            lcout => chessboardpixel_un152_pixel_24,
            ltout => OPEN,
            carryin => un5_visiblex_cry_2,
            carryout => un5_visiblex_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10453\,
            in3 => \N__10417\,
            lcout => charx_if_generate_plus_mult1_un54_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_3,
            carryout => un5_visiblex_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10410\,
            in3 => \N__10372\,
            lcout => charx_if_generate_plus_mult1_un47_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_4,
            carryout => un5_visiblex_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16395\,
            in2 => \N__10369\,
            in3 => \N__10333\,
            lcout => charx_if_generate_plus_mult1_un40_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_5,
            carryout => un5_visiblex_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10311\,
            in2 => \_gnd_net_\,
            in3 => \N__10285\,
            lcout => charx_if_generate_plus_mult1_un33_sum,
            ltout => OPEN,
            carryin => un5_visiblex_cry_6,
            carryout => un5_visiblex_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16396\,
            in2 => \N__10282\,
            in3 => \N__10249\,
            lcout => charx_if_generate_plus_mult1_un26_sum,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => un5_visiblex_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10735\,
            in2 => \_gnd_net_\,
            in3 => \N__10714\,
            lcout => \CO3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_5_c_RNIR332_1_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13876\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_3_bm_2_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13417\,
            in2 => \N__16030\,
            in3 => \N__14750\,
            lcout => OPEN,
            ltout => \un116_pixel_3_bm_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_3_ns_2_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14949\,
            in2 => \N__10711\,
            in3 => \N__11662\,
            lcout => un116_pixel_3_ns_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111001010000"
        )
    port map (
            in0 => \N__15814\,
            in1 => \N__10696\,
            in2 => \N__10708\,
            in3 => \N__15355\,
            lcout => \N_345_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_16_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101010011"
        )
    port map (
            in0 => \N__15354\,
            in1 => \N__15813\,
            in2 => \N__14995\,
            in3 => \N__15585\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un116_pixel_4_ns_1_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_12_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101010101110"
        )
    port map (
            in0 => \N__14950\,
            in1 => \N__14255\,
            in2 => \N__10699\,
            in3 => \N__16029\,
            lcout => \N_347_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g2_1_0_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__15592\,
            in1 => \N__16024\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \un114_pixel_1_0_3__g2_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJPPPPD1_0_3_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010001000010"
        )
    port map (
            in0 => \N__12264\,
            in1 => \N__12281\,
            in2 => \N__10686\,
            in3 => \N__10669\,
            lcout => OPEN,
            ltout => \font_un28_pixel_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_i_m2_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101100101000"
        )
    port map (
            in0 => \N__10780\,
            in1 => \N__14954\,
            in2 => \N__10774\,
            in3 => \N__14269\,
            lcout => \N_346_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_5_am_6_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011111111100"
        )
    port map (
            in0 => \N__15591\,
            in1 => \N__15337\,
            in2 => \N__15816\,
            in3 => \N__16019\,
            lcout => OPEN,
            ltout => \un116_pixel_5_am_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_5_ns_6_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14753\,
            in2 => \N__10771\,
            in3 => \N__11812\,
            lcout => \N_379\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_0_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100101000"
        )
    port map (
            in0 => \N__12280\,
            in1 => \N__10768\,
            in2 => \N__10762\,
            in3 => \N__12263\,
            lcout => font_un28_pixel_0_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_2_ns_1_2_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101111100"
        )
    port map (
            in0 => \N__15590\,
            in1 => \N__15336\,
            in2 => \N__15815\,
            in3 => \N__16017\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un116_pixel_2_ns_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_2_ns_2_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__16018\,
            in1 => \N__14752\,
            in2 => \N__10753\,
            in3 => \N__13418\,
            lcout => \N_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_5_ns_1_2_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__14741\,
            in1 => \N__15580\,
            in2 => \_gnd_net_\,
            in3 => \N__15334\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un116_pixel_5_ns_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_5_ns_2_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001101000000"
        )
    port map (
            in0 => \N__16021\,
            in1 => \N__14742\,
            in2 => \N__10750\,
            in3 => \N__15812\,
            lcout => un116_pixel_5_ns_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_5_ns_1_4_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100000111100"
        )
    port map (
            in0 => \N__15586\,
            in1 => \N__15335\,
            in2 => \N__15817\,
            in3 => \N__16022\,
            lcout => OPEN,
            ltout => \un116_pixel_5_ns_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI2L0T663_0_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000110101001"
        )
    port map (
            in0 => \N__16023\,
            in1 => \N__14743\,
            in2 => \N__10840\,
            in3 => \N__13422\,
            lcout => \beamY_RNI2L0T663Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIPU5VF83_1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010011"
        )
    port map (
            in0 => \N__10837\,
            in1 => \N__10831\,
            in2 => \N__15012\,
            in3 => \N__13292\,
            lcout => OPEN,
            ltout => \un116_pixel_7_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIVU1O9R_1_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__13293\,
            in1 => \N__10786\,
            in2 => \N__10825\,
            in3 => \N__10822\,
            lcout => \beamY_RNIVU1O9RZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI57H3N31_0_1_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__14901\,
            in1 => \N__11793\,
            in2 => \N__13306\,
            in3 => \N__10804\,
            lcout => OPEN,
            ltout => \beamY_RNI57H3N31_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1J75181_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10816\,
            in2 => \N__10807\,
            in3 => \N__10795\,
            lcout => \beamY_RNI1J75181Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI896FQ3_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__14217\,
            in1 => \N__11938\,
            in2 => \N__14759\,
            in3 => \N__11074\,
            lcout => \beamY_RNI896FQ3Z0Z_0\,
            ltout => \beamY_RNI896FQ3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI57H3N31_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011111111"
        )
    port map (
            in0 => \N__11794\,
            in1 => \N__14900\,
            in2 => \N__10798\,
            in3 => \N__13295\,
            lcout => \beamY_RNI57H3N31Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIAK9BMC1_0_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110011001"
        )
    port map (
            in0 => \N__15754\,
            in1 => \N__14630\,
            in2 => \_gnd_net_\,
            in3 => \N__15584\,
            lcout => OPEN,
            ltout => \un116_pixel_2_ns_1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIGO5PPV_0_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000111010"
        )
    port map (
            in0 => \N__15296\,
            in1 => \N__15755\,
            in2 => \N__10789\,
            in3 => \N__13363\,
            lcout => \beamY_RNIGO5PPVZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un114_pixel_3_i_m2_i_m2_6_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110101100110"
        )
    port map (
            in0 => \N__15753\,
            in1 => \N__15295\,
            in2 => \N__14244\,
            in3 => \N__16020\,
            lcout => \N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_1_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001101100"
        )
    port map (
            in0 => \N__11026\,
            in1 => \N__14902\,
            in2 => \N__14702\,
            in3 => \N__10977\,
            lcout => \beamYZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11882\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_1_c_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13599\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_2_s_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11139\,
            in2 => \N__10900\,
            in3 => \N__10912\,
            lcout => if_generate_plus_mult1_un68_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_cry_3_s_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11125\,
            in2 => \N__15544\,
            in3 => \N__10909\,
            lcout => if_generate_plus_mult1_un68_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_5_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15249\,
            in1 => \N__11140\,
            in2 => \N__11116\,
            in3 => \N__10906\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_s_5_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11104\,
            in2 => \_gnd_net_\,
            in3 => \N__10903\,
            lcout => un5_rowlto2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_i_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11538\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_row_8_7_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110000"
        )
    port map (
            in0 => \N__15287\,
            in1 => \N__10890\,
            in2 => \N__15545\,
            in3 => \N__16016\,
            lcout => \un114_pixel_1_0_3__un4_row_8_7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_rowlto3_sbtinv_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15492\,
            lcout => un5_rowlto3_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11537\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_8_0_\,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_2_s_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11131\,
            in2 => \N__11092\,
            in3 => \N__11119\,
            lcout => if_generate_plus_mult1_un61_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_cry_3_s_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11353\,
            in2 => \N__12508\,
            in3 => \N__11107\,
            lcout => if_generate_plus_mult1_un61_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_axb_5_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15499\,
            in1 => \N__11091\,
            in2 => \N__11338\,
            in3 => \N__11098\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_s_5_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11320\,
            in2 => \_gnd_net_\,
            in3 => \N__11095\,
            lcout => un5_rowlto3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12503\,
            lcout => column_1_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__N_37_i_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__15081\,
            in1 => \N__14030\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_37_i\,
            ltout => OPEN,
            carryin => \bfn_7_9_0_\,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57K_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11290\,
            in2 => \N__11211\,
            in3 => \N__11077\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_1_c_RNIU57KZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15Q_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11257\,
            in2 => \N__11230\,
            in3 => \N__11251\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_2_c_RNIG15QZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8BLE3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11193\,
            in1 => \N__11248\,
            in2 => \N__11212\,
            in3 => \N__11242\,
            lcout => charx_if_generate_plus_mult1_un40_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un33_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un33_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11239\,
            in2 => \_gnd_net_\,
            in3 => \N__11233\,
            lcout => \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNIZ0Z65072\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un26_sum_cry_4_c_RNIISU5_0_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11225\,
            lcout => charx_if_generate_plus_mult1_un26_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un33_sum_cry_4_c_RNI65072_0_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11192\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13858\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_10_0_\,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEB2_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11296\,
            in2 => \N__11157\,
            in3 => \N__11197\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_1_c_RNIEKEBZ0Z2\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLIT2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11194\,
            in2 => \N__11176\,
            in3 => \N__11167\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_2_c_RNIGLITZ0Z2\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_3_c_RNIPCKK6_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11456\,
            in1 => \N__11164\,
            in2 => \N__11158\,
            in3 => \N__11143\,
            lcout => charx_if_generate_plus_mult1_un47_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un40_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un40_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11305\,
            in2 => \_gnd_net_\,
            in3 => \N__11299\,
            lcout => \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2HZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14031\,
            lcout => charx_if_generate_plus_mult1_un33_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15065\,
            lcout => charx_if_generate_plus_mult1_un26_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__12896\,
            in1 => \N__14032\,
            in2 => \_gnd_net_\,
            in3 => \N__16153\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_1_c_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13868\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11284\,
            in2 => \N__11380\,
            in3 => \N__11278\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_2,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_1,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12832\,
            in2 => \N__11371\,
            in3 => \N__11275\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_3,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_2,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11272\,
            in2 => \N__11362\,
            in3 => \N__11263\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_4,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_0_cry_3,
            carryout => column_1_if_generate_plus_mult1_un47_sum_0_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_s_5_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16152\,
            in2 => \_gnd_net_\,
            in3 => \N__11260\,
            lcout => column_1_if_generate_plus_mult1_un47_sum0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_2_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14038\,
            lcout => un5_visiblex_i_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__16138\,
            in1 => \N__12924\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => if_generate_plus_mult1_un47_sum_0_cry_3_ma,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__16151\,
            in1 => \N__15077\,
            in2 => \N__12935\,
            in3 => \N__14039\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11652\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13033\,
            in2 => \N__12963\,
            in3 => \N__11341\,
            lcout => if_generate_plus_mult1_un54_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13005\,
            in2 => \N__12991\,
            in3 => \N__11323\,
            lcout => if_generate_plus_mult1_un54_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12499\,
            in1 => \N__11476\,
            in2 => \N__12964\,
            in3 => \N__11311\,
            lcout => \column_1_if_generate_plus_mult1_un61_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13018\,
            in2 => \_gnd_net_\,
            in3 => \N__11308\,
            lcout => if_generate_plus_mult1_un54_sum_s_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un40_sum_cry_4_c_RNIMP2H3_0_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11457\,
            lcout => charx_if_generate_plus_mult1_un40_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_4_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100111000011"
        )
    port map (
            in0 => \N__11485\,
            in1 => \N__13004\,
            in2 => \N__14134\,
            in3 => \N__16154\,
            lcout => OPEN,
            ltout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11479\,
            in3 => \N__12956\,
            lcout => if_generate_plus_mult1_un54_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11650\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0O3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11470\,
            in2 => \N__11412\,
            in3 => \N__11461\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_1_c_RNI3Q0OZ0Z3\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCD16_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11458\,
            in2 => \N__11437\,
            in3 => \N__11425\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_2_c_RNINCDZ0Z16\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_3_c_RNI8V4DD_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11604\,
            in1 => \N__11422\,
            in2 => \N__11413\,
            in3 => \N__11398\,
            lcout => charx_if_generate_plus_mult1_un54_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un47_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11395\,
            in2 => \_gnd_net_\,
            in3 => \N__11386\,
            lcout => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6\,
            ltout => \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIPZ0Z6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un47_sum_cry_4_c_RNIEFIP6_0_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11383\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_4_c_RNIP022_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11651\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11545\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLM67_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11614\,
            in2 => \N__11574\,
            in3 => \N__11608\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_1_c_RNINLMZ0Z67\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSA_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11605\,
            in2 => \N__11593\,
            in3 => \N__11584\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_2_c_RNI2HMSAZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_3_c_RNIIGEUQ_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11700\,
            in1 => \N__11581\,
            in2 => \N__11575\,
            in3 => \N__11560\,
            lcout => charx_if_generate_plus_mult1_un61_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un54_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11557\,
            in2 => \_gnd_net_\,
            in3 => \N__11551\,
            lcout => \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAODZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_3_c_RNINT02_0_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11546\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13603\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRD_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11494\,
            in2 => \N__11682\,
            in3 => \N__11488\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_1_c_RNI0NKRDZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0L_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11731\,
            in2 => \N__11701\,
            in3 => \N__11725\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_2_c_RNI1HB0LZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_3_c_RNIGJ7MJ1_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13161\,
            in1 => \N__11722\,
            in2 => \N__11683\,
            in3 => \N__11716\,
            lcout => charx_if_generate_plus_mult1_un68_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un61_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11713\,
            in2 => \_gnd_net_\,
            in3 => \N__11707\,
            lcout => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0\,
            ltout => \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un61_sum_cry_4_c_RNI35RVQ_0_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11704\,
            in3 => \_gnd_net_\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un54_sum_cry_4_c_RNIRAAOD_0_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11696\,
            lcout => charx_if_generate_plus_mult1_un54_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VSyncZ0_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12060\,
            lcout => \VSync_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11884\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_3_am_2_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011100001"
        )
    port map (
            in0 => \N__15808\,
            in1 => \N__15382\,
            in2 => \N__14776\,
            in3 => \N__16028\,
            lcout => un116_pixel_3_am_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_2_0_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001101100"
        )
    port map (
            in0 => \N__13424\,
            in1 => \N__14757\,
            in2 => \N__15015\,
            in3 => \N__13228\,
            lcout => \N_368_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_13_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__16012\,
            in1 => \N__13045\,
            in2 => \N__14777\,
            in3 => \N__13423\,
            lcout => OPEN,
            ltout => \N_1556_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_11_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__15003\,
            in1 => \N__14278\,
            in2 => \N__11782\,
            in3 => \_gnd_net_\,
            lcout => \N_389_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_0_0_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110101"
        )
    port map (
            in0 => \N__11779\,
            in1 => \N__13213\,
            in2 => \N__11770\,
            in3 => \N__13303\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__font_un126_pixel_1_d_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__13304\,
            in1 => \N__11761\,
            in2 => \N__11755\,
            in3 => \N__11752\,
            lcout => OPEN,
            ltout => \g0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_i_m2_0_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__14758\,
            in1 => \N__11746\,
            in2 => \N__11740\,
            in3 => \N__13305\,
            lcout => \N_400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__m18_0_m2_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101101010101"
        )
    port map (
            in0 => \N__15791\,
            in1 => \N__15589\,
            in2 => \_gnd_net_\,
            in3 => \N__15333\,
            lcout => \N_36\,
            ltout => \N_36_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_1_4_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011001110"
        )
    port map (
            in0 => \N__16011\,
            in1 => \N__14751\,
            in2 => \N__11737\,
            in3 => \N__13234\,
            lcout => un116_pixel_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIC1MEAP2_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__14461\,
            in1 => \_gnd_net_\,
            in2 => \N__13426\,
            in3 => \N__14800\,
            lcout => OPEN,
            ltout => \un116_pixel_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNILBST4T2_1_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__14986\,
            in1 => \N__13432\,
            in2 => \N__11734\,
            in3 => \N__11806\,
            lcout => \beamY_RNILBST4T2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__N_315_i_i_a3_0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15577\,
            in2 => \_gnd_net_\,
            in3 => \N__15326\,
            lcout => \N_563\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010111110000"
        )
    port map (
            in0 => \N__13543\,
            in1 => \_gnd_net_\,
            in2 => \N__13513\,
            in3 => \N__13464\,
            lcout => font_un3_pixel_29,
            ltout => \font_un3_pixel_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_7_x1_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101001111"
        )
    port map (
            in0 => \N__13318\,
            in1 => \N__14987\,
            in2 => \N__11815\,
            in3 => \N__13334\,
            lcout => un116_pixel_7_x1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_5_bm_6_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001110010111110"
        )
    port map (
            in0 => \N__16000\,
            in1 => \N__15807\,
            in2 => \N__15384\,
            in3 => \N__14238\,
            lcout => un116_pixel_5_bm_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__m5_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15578\,
            in2 => \_gnd_net_\,
            in3 => \N__15998\,
            lcout => \N_325\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_4_bm_1_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011011110110"
        )
    port map (
            in0 => \N__15999\,
            in1 => \N__15806\,
            in2 => \N__15383\,
            in3 => \N__15579\,
            lcout => un116_pixel_4_bm_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI1C50FS3_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011111010"
        )
    port map (
            in0 => \N__13381\,
            in1 => \N__13375\,
            in2 => \N__14775\,
            in3 => \N__14161\,
            lcout => OPEN,
            ltout => \beamY_RNI1C50FS3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un126_pixel_2_bm_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13204\,
            in2 => \N__11800\,
            in3 => \N__13300\,
            lcout => font_un126_pixel_2_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIG8FT9A2_0_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100000101"
        )
    port map (
            in0 => \N__15770\,
            in1 => \N__15588\,
            in2 => \N__14774\,
            in3 => \N__15288\,
            lcout => OPEN,
            ltout => \un116_pixel_3_bm_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIOHI2NG_0_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101110100"
        )
    port map (
            in0 => \N__16009\,
            in1 => \N__14736\,
            in2 => \N__11797\,
            in3 => \N__15294\,
            lcout => \beamY_RNIOHI2NGZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_2_ns_0_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14737\,
            in1 => \N__13624\,
            in2 => \_gnd_net_\,
            in3 => \N__15442\,
            lcout => OPEN,
            ltout => \N_364_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI57H3N31_1_1_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__14903\,
            in1 => \N__13369\,
            in2 => \N__11950\,
            in3 => \N__13299\,
            lcout => OPEN,
            ltout => \un116_pixel_7_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI7OE17C_0_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__13301\,
            in1 => \N__14545\,
            in2 => \N__11947\,
            in3 => \N__11944\,
            lcout => \beamY_RNI7OE17CZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__column_0111_1_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__16010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15769\,
            lcout => column_0111_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un126_pixel_6_am_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110101001000"
        )
    port map (
            in0 => \N__13541\,
            in1 => \N__13240\,
            in2 => \N__13465\,
            in3 => \N__11932\,
            lcout => OPEN,
            ltout => \font_un126_pixel_6_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_1_1_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100010"
        )
    port map (
            in0 => \N__12023\,
            in1 => \N__11821\,
            in2 => \N__11926\,
            in3 => \N__12127\,
            lcout => OPEN,
            ltout => \N_1075_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_4_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__11923\,
            in1 => \N__12310\,
            in2 => \N__11911\,
            in3 => \N__12067\,
            lcout => OPEN,
            ltout => \Pixel_r_rn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PixelZ0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11908\,
            in2 => \N__11899\,
            in3 => \N__12031\,
            lcout => \Pixel_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_7_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010101110101"
        )
    port map (
            in0 => \N__11839\,
            in1 => \N__11827\,
            in2 => \N__12025\,
            in3 => \N__13186\,
            lcout => \un114_pixel_1_0_3__font_un126_pixel_7_d_ns_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNI90K6F01_2_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12292\,
            in2 => \_gnd_net_\,
            in3 => \N__12265\,
            lcout => chary_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un126_pixel_6_bm_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__13540\,
            in1 => \N__13460\,
            in2 => \N__12145\,
            in3 => \N__12136\,
            lcout => font_un126_pixel_6_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIAV9A43_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14451\,
            in2 => \_gnd_net_\,
            in3 => \N__13663\,
            lcout => charx_if_generate_plus_mult1_un1_sum_axb1,
            ltout => \charx_if_generate_plus_mult1_un1_sum_axb1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNIEUFG5F_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13509\,
            in2 => \N__12121\,
            in3 => \N__13458\,
            lcout => OPEN,
            ltout => \r_i1_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un126_pixel_m_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110001001100"
        )
    port map (
            in0 => \N__13492\,
            in1 => \N__12117\,
            in2 => \N__12094\,
            in3 => \N__12018\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un126_pixel_m_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__12360\,
            in1 => \N__12342\,
            in2 => \N__12091\,
            in3 => \N__12370\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__font_un126_pixel_m_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un126_pixel_m_3_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000001100000"
        )
    port map (
            in0 => \N__14974\,
            in1 => \N__12088\,
            in2 => \N__12076\,
            in3 => \N__12073\,
            lcout => \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3\,
            ltout => \un114_pixel_1_0_3__font_un126_pixel_mZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Pixel_RNO_0_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__12061\,
            in1 => \N__12306\,
            in2 => \N__12034\,
            in3 => \N__12826\,
            lcout => \Pixel_r_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un57_pixel_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__13459\,
            in1 => \N__13542\,
            in2 => \_gnd_net_\,
            in3 => \N__12019\,
            lcout => \un114_pixel_1_0_3__font_un57_pixelZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_row_8_3_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000001010000"
        )
    port map (
            in0 => \N__12601\,
            in1 => \N__12820\,
            in2 => \N__12478\,
            in3 => \N__12691\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un4_row_8Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_row_8_7_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12730\,
            in1 => \N__12447\,
            in2 => \N__12703\,
            in3 => \N__12700\,
            lcout => \un114_pixel_1_0_3__un4_row_8Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_row_8_2_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__12690\,
            in1 => \N__12600\,
            in2 => \N__12853\,
            in3 => \N__12507\,
            lcout => \un114_pixel_1_0_3__un4_row_8Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_row_8_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100100000000"
        )
    port map (
            in0 => \N__12469\,
            in1 => \N__12448\,
            in2 => \N__12418\,
            in3 => \N__12376\,
            lcout => \un114_pixel_1_0_3__un4_rowZ0Z_8\,
            ltout => \un114_pixel_1_0_3__un4_rowZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__Pixel_3_sqmuxa_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111100000000"
        )
    port map (
            in0 => \N__12364\,
            in1 => \N__12343\,
            in2 => \N__12322\,
            in3 => \N__12319\,
            lcout => \Pixel_3_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_1_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101111110000"
        )
    port map (
            in0 => \N__14450\,
            in1 => \N__13719\,
            in2 => \N__13690\,
            in3 => \N__13659\,
            lcout => font_un3_pixel_if_generate_plus_mult1_un25_sum_s_4_sf,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14425\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_10_0_\,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46K1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12859\,
            in2 => \N__12841\,
            in3 => \N__12295\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIEV46KZ0Z1\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9F2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13177\,
            in2 => \N__13081\,
            in3 => \N__12877\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI9CS9FZ0Z2\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_inv_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13141\,
            in2 => \N__12874\,
            in3 => \N__13077\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_invZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPAC843_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13105\,
            in2 => \_gnd_net_\,
            in3 => \N__12865\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843\,
            ltout => \charx_if_generate_plus_mult1_un75_sum_cry_4_c_RNIPACZ0Z843_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNO_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111101010000"
        )
    port map (
            in0 => \N__14426\,
            in1 => \_gnd_net_\,
            in2 => \N__12862\,
            in3 => \N__13713\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_1_c_RNIJNU1_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15148\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_N_858_i_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16184\,
            lcout => \N_858_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un4_row_8_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__16186\,
            in1 => \N__12923\,
            in2 => \N__14098\,
            in3 => \N__12982\,
            lcout => \un114_pixel_1_0_3__un4_row_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13076\,
            lcout => charx_if_generate_plus_mult1_un68_sum_i_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011111010"
        )
    port map (
            in0 => \N__14004\,
            in1 => \N__12919\,
            in2 => \N__12934\,
            in3 => \N__16185\,
            lcout => if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111101110"
        )
    port map (
            in0 => \N__14003\,
            in1 => \N__12918\,
            in2 => \_gnd_net_\,
            in3 => \N__16183\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_3_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_2_sx_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100001001"
        )
    port map (
            in0 => \N__13886\,
            in1 => \N__14089\,
            in2 => \N__16209\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \column_1_if_generate_plus_mult1_un54_sum_axb_2_sxZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_2_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001101"
        )
    port map (
            in0 => \N__16201\,
            in1 => \N__13887\,
            in2 => \N__13039\,
            in3 => \N__12981\,
            lcout => OPEN,
            ltout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13036\,
            in3 => \N__12955\,
            lcout => if_generate_plus_mult1_un54_sum_axb_2_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_m_5_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16191\,
            in2 => \N__14097\,
            in3 => \N__12979\,
            lcout => if_generate_plus_mult1_un47_sum_m_5,
            ltout => \if_generate_plus_mult1_un47_sum_m_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_5_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110100101"
        )
    port map (
            in0 => \N__14110\,
            in1 => \N__13027\,
            in2 => \N__13021\,
            in3 => \N__16203\,
            lcout => \column_1_if_generate_plus_mult1_un54_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__16202\,
            in1 => \N__13012\,
            in2 => \N__13819\,
            in3 => \N__13006\,
            lcout => if_generate_plus_mult1_un54_sum_axb_3_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_N_584_i_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101010011"
        )
    port map (
            in0 => \N__12980\,
            in1 => \N__14093\,
            in2 => \N__16208\,
            in3 => \_gnd_net_\,
            lcout => \N_584_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16190\,
            in2 => \N__14005\,
            in3 => \N__12936\,
            lcout => if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15155\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5R_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13051\,
            in2 => \N__13119\,
            in3 => \N__13165\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_1_c_RNID2L5RZ0\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_1,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BV81_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13162\,
            in2 => \N__13150\,
            in3 => \N__13129\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_2_c_RNIP0BVZ0Z81\,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_2,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_3_c_RNI3P7U33_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13070\,
            in1 => \N__13126\,
            in2 => \N__13120\,
            in3 => \N__13093\,
            lcout => charx_if_generate_plus_mult1_un75_sum_axb_5,
            ltout => OPEN,
            carryin => charx_if_generate_plus_mult1_un68_sum_cry_3,
            carryout => charx_if_generate_plus_mult1_un68_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJ1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13090\,
            in2 => \_gnd_net_\,
            in3 => \N__13084\,
            lcout => \charx_if_generate_plus_mult1_un68_sum_cry_4_c_RNI8S4QJZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_2_c_RNILQV1_0_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13611\,
            lcout => charx_if_generate_plus_mult1_un61_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_i_m2_1_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101110010"
        )
    port map (
            in0 => \N__16002\,
            in1 => \N__14239\,
            in2 => \N__15405\,
            in3 => \N__15793\,
            lcout => \N_41_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g1_4_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__15795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15608\,
            lcout => \un114_pixel_1_0_3__g1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__column_0111_0_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15792\,
            in1 => \N__15385\,
            in2 => \_gnd_net_\,
            in3 => \N__16001\,
            lcout => column_0111_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_3_1_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011110001"
        )
    port map (
            in0 => \N__15796\,
            in1 => \N__15389\,
            in2 => \N__15014\,
            in3 => \N__16003\,
            lcout => un116_pixel_3_ns_1_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_17_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111101110010"
        )
    port map (
            in0 => \N__16004\,
            in1 => \N__14240\,
            in2 => \N__15406\,
            in3 => \N__15794\,
            lcout => OPEN,
            ltout => \N_1583_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_14_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__14999\,
            in1 => \N__13222\,
            in2 => \N__13216\,
            in3 => \N__15393\,
            lcout => \N_26_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_2_am_1_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101000100"
        )
    port map (
            in0 => \N__15395\,
            in1 => \N__15804\,
            in2 => \N__14254\,
            in3 => \N__16007\,
            lcout => OPEN,
            ltout => \un116_pixel_2_amZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_6_1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100111001000"
        )
    port map (
            in0 => \N__14985\,
            in1 => \N__13345\,
            in2 => \N__13207\,
            in3 => \N__13351\,
            lcout => un116_pixel_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_4_0_15__m15_0_a3_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14237\,
            in1 => \N__15805\,
            in2 => \_gnd_net_\,
            in3 => \N__16008\,
            lcout => OPEN,
            ltout => \column_0001_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIT81CMJ2_1_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110100010"
        )
    port map (
            in0 => \N__14984\,
            in1 => \N__14746\,
            in2 => \N__13198\,
            in3 => \N__13335\,
            lcout => OPEN,
            ltout => \beamY_RNIT81CMJ2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__font_un126_pixel_2_am_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13195\,
            in2 => \N__13189\,
            in3 => \N__13294\,
            lcout => font_un126_pixel_2_am,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_4_am_1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000110111011"
        )
    port map (
            in0 => \N__15394\,
            in1 => \N__15803\,
            in2 => \N__14253\,
            in3 => \N__16005\,
            lcout => un116_pixel_4_am_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__m20_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__16006\,
            in1 => \N__14745\,
            in2 => \_gnd_net_\,
            in3 => \N__13425\,
            lcout => \N_374_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_5_am_5_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010001000"
        )
    port map (
            in0 => \N__16014\,
            in1 => \N__14221\,
            in2 => \N__15404\,
            in3 => \N__15757\,
            lcout => \un116_pixel_5_amZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_2_am_5_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__15758\,
            in1 => \N__16015\,
            in2 => \N__14246\,
            in3 => \N__15380\,
            lcout => \un116_pixel_2_amZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_5_ns_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111000000"
        )
    port map (
            in0 => \N__15381\,
            in1 => \N__13618\,
            in2 => \N__14773\,
            in3 => \N__15760\,
            lcout => \N_385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_2_bm_1_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__15759\,
            in1 => \N__13362\,
            in2 => \_gnd_net_\,
            in3 => \N__15375\,
            lcout => \un116_pixel_2_bmZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_6_1_1_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110000101"
        )
    port map (
            in0 => \N__14729\,
            in1 => \N__13552\,
            in2 => \N__14975\,
            in3 => \N__15761\,
            lcout => \un114_pixel_1_0_3__un116_pixel_6_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_7_x0_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000000000"
        )
    port map (
            in0 => \N__13339\,
            in1 => \N__13317\,
            in2 => \N__14976\,
            in3 => \N__13302\,
            lcout => OPEN,
            ltout => \un116_pixel_7_x0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_7_ns_0_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14473\,
            in2 => \N__13249\,
            in3 => \N__13246\,
            lcout => un116_pixel_7_ns_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_2_bm_0_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011100110"
        )
    port map (
            in0 => \N__15756\,
            in1 => \N__16013\,
            in2 => \N__14245\,
            in3 => \N__15376\,
            lcout => un116_pixel_2_bm_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_5_ns_1_0_0_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001111010011"
        )
    port map (
            in0 => \N__15594\,
            in1 => \N__15919\,
            in2 => \N__14744\,
            in3 => \N__15302\,
            lcout => \un114_pixel_1_0_3__un116_pixel_5_ns_1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un68_sum_i_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13607\,
            lcout => \column_1_if_generate_plus_mult1_un68_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_6_1_1_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__15593\,
            in1 => \N__15918\,
            in2 => \_gnd_net_\,
            in3 => \N__15301\,
            lcout => \un114_pixel_1_0_3__un116_pixel_6_1_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13536\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSO4_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13749\,
            in2 => \N__13729\,
            in3 => \N__13495\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1_c_RNI1JJSOZ0Z4\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3E987_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13798\,
            in2 => \N__13482\,
            in3 => \N__13486\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2_c_RNIV3EZ0Z987\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNIN803_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13750\,
            in2 => \N__13789\,
            in3 => \N__13748\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_c_RNINZ0Z803\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CI987_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13776\,
            in1 => \N__13762\,
            in2 => \N__13483\,
            in3 => \N__13468\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNI3CIZ0Z987\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13807\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8T77_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13633\,
            in3 => \N__13792\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1_c_RNILD8TZ0Z77\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_1,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNO_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16397\,
            in2 => \N__13738\,
            in3 => \N__13780\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un32_sum_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_2,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_LUT4_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13777\,
            in3 => \N__13756\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_3,
            carryout => font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_LUT4_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13753\,
            lcout => \font_un3_pixel_if_generate_plus_mult1_un25_sum_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000001111"
        )
    port map (
            in0 => \N__14445\,
            in1 => \N__13715\,
            in2 => \N__13689\,
            in3 => \N__13657\,
            lcout => \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_1_c_RNIOUEGO4_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110100101"
        )
    port map (
            in0 => \N__13658\,
            in1 => \_gnd_net_\,
            in2 => \N__13720\,
            in3 => \N__14446\,
            lcout => charx_i_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \charx_if_generate_plus_mult1_un75_sum_cry_2_c_RNI1BBQ77_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011010000001111"
        )
    port map (
            in0 => \N__14444\,
            in1 => \N__13714\,
            in2 => \N__13688\,
            in3 => \N__13656\,
            lcout => charx_i_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13888\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_11_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUH2_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13894\,
            in2 => \N__14073\,
            in3 => \N__13948\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNI9CUHZ0Z2\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIV6153_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14365\,
            in2 => \N__13984\,
            in3 => \N__13933\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIVZ0Z6153\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNISAMG7_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__13910\,
            in1 => \N__13969\,
            in2 => \N__14074\,
            in3 => \N__13921\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un68_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6T3_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14380\,
            in2 => \_gnd_net_\,
            in3 => \N__13918\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNIGP6TZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_3_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14057\,
            lcout => un5_visiblex_i_0_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_6_c_RNIT642_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14058\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13885\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_2_s_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16198\,
            in2 => \N__13828\,
            in3 => \N__13810\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_2,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_1,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14149\,
            in2 => \N__14143\,
            in3 => \N__14122\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_3,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_2,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16199\,
            in2 => \N__14119\,
            in3 => \N__14104\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_4,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un47_sum_1_cry_3,
            carryout => column_1_if_generate_plus_mult1_un47_sum_1_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un47_sum_1_s_5_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000001111111"
        )
    port map (
            in0 => \N__16200\,
            in1 => \N__14059\,
            in2 => \N__15106\,
            in3 => \N__14101\,
            lcout => column_1_if_generate_plus_mult1_un47_sum1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_0_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14360\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_0_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16236\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__SUM4_3_i_a2_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14048\,
            in2 => \_gnd_net_\,
            in3 => \N__15097\,
            lcout => \N_66\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5L_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14388\,
            in2 => \N__14344\,
            in3 => \N__13972\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIIV5LZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7J31_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16240\,
            in2 => \N__16429\,
            in3 => \N__13960\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIU7JZ0Z31\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI8U9I3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__14361\,
            in1 => \N__14389\,
            in2 => \N__16276\,
            in3 => \N__14371\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un61_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7G052_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16258\,
            in2 => \_gnd_net_\,
            in3 => \N__14368\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI7GZ0Z052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_7_c_RNIV952_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15098\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_Clock12MHz_c_g_THRU_LUT4_0_LC_11_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14335\,
            lcout => \GB_BUFFER_Clock12MHz_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_15_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000011001"
        )
    port map (
            in0 => \N__15402\,
            in1 => \N__15789\,
            in2 => \N__14779\,
            in3 => \N__15996\,
            lcout => \N_1557_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIKBQK731_0_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__14769\,
            in1 => \N__15616\,
            in2 => \_gnd_net_\,
            in3 => \N__15401\,
            lcout => un116_pixel_2_ns_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__g0_i_m2_2_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101101100110"
        )
    port map (
            in0 => \N__15403\,
            in1 => \N__15790\,
            in2 => \N__14260\,
            in3 => \N__15997\,
            lcout => \N_41_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_5_bm_5_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000000000"
        )
    port map (
            in0 => \N__15397\,
            in1 => \N__15693\,
            in2 => \N__14256\,
            in3 => \N__15982\,
            lcout => OPEN,
            ltout => \un116_pixel_5_bmZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJEPU0R2_1_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100101011101"
        )
    port map (
            in0 => \N__15010\,
            in1 => \N__14766\,
            in2 => \N__14164\,
            in3 => \N__14491\,
            lcout => un116_pixel_6_ns_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__m33_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010000010001"
        )
    port map (
            in0 => \N__15398\,
            in1 => \N__15695\,
            in2 => \N__15618\,
            in3 => \N__15983\,
            lcout => \un114_pixel_6_1_5__N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_2_bm_5_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__15692\,
            in1 => \N__15609\,
            in2 => \_gnd_net_\,
            in3 => \N__15396\,
            lcout => \un116_pixel_2_bmZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__m24_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010011001"
        )
    port map (
            in0 => \N__15399\,
            in1 => \N__15694\,
            in2 => \N__15619\,
            in3 => \N__15984\,
            lcout => OPEN,
            ltout => \un114_pixel_7_1_7__N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_3_ns_1_0_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000011101"
        )
    port map (
            in0 => \N__15696\,
            in1 => \N__14767\,
            in2 => \N__14485\,
            in3 => \N__15400\,
            lcout => OPEN,
            ltout => \un114_pixel_1_0_3__un116_pixel_3_ns_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_3_ns_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001011011011"
        )
    port map (
            in0 => \N__14768\,
            in1 => \N__15011\,
            in2 => \N__14482\,
            in3 => \N__14479\,
            lcout => \N_371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIJUCG3J3_1_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001100110"
        )
    port map (
            in0 => \N__15009\,
            in1 => \N__14765\,
            in2 => \_gnd_net_\,
            in3 => \N__15022\,
            lcout => \beamY_RNIJUCG3J3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_1_c_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14452\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14395\,
            in2 => \N__15121\,
            in3 => \N__15861\,
            lcout => \G_345\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_3_c_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14524\,
            in2 => \N__15917\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15034\,
            in2 => \N__14503\,
            in3 => \N__15862\,
            lcout => \G_346\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un82_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un82_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_s_5_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16051\,
            in2 => \_gnd_net_\,
            in3 => \N__15028\,
            lcout => un5_rowlto0,
            ltout => \un5_rowlto0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un116_pixel_1_bm_1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011000011"
        )
    port map (
            in0 => \N__15587\,
            in1 => \N__15356\,
            in2 => \N__15025\,
            in3 => \N__15866\,
            lcout => \un116_pixel_1_bmZ0Z_1\,
            ltout => \un116_pixel_1_bmZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIV622TR_1_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111101110"
        )
    port map (
            in0 => \N__15867\,
            in1 => \N__14920\,
            in2 => \N__14803\,
            in3 => \N__14761\,
            lcout => \beamY_RNIV622TRZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \beamY_RNIITCG3J3_0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000111010000"
        )
    port map (
            in0 => \N__15728\,
            in1 => \N__14788\,
            in2 => \N__14778\,
            in3 => \N__15868\,
            lcout => \beamY_RNIITCG3J3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_1_c_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15162\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_2_s_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15169\,
            in2 => \N__14536\,
            in3 => \N__14518\,
            lcout => if_generate_plus_mult1_un75_sum_cry_2_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_1,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_cry_3_s_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15300\,
            in2 => \N__14515\,
            in3 => \N__14494\,
            lcout => if_generate_plus_mult1_un75_sum_cry_3_s,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_2,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un82_sum_axb_5_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__15869\,
            in1 => \N__15412\,
            in2 => \N__15430\,
            in3 => \N__16045\,
            lcout => \column_1_if_generate_plus_mult1_un82_sum_axbZ0Z_5\,
            ltout => OPEN,
            carryin => column_1_if_generate_plus_mult1_un75_sum_cry_3,
            carryout => column_1_if_generate_plus_mult1_un75_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_s_5_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16042\,
            in2 => \_gnd_net_\,
            in3 => \N__16033\,
            lcout => un5_rowlto1,
            ltout => \un5_rowlto1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un114_pixel_1_0_3__un116_pixel_2_am_0_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011011110"
        )
    port map (
            in0 => \N__15684\,
            in1 => \N__15299\,
            in2 => \N__15622\,
            in3 => \N__15617\,
            lcout => un116_pixel_2_am_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_axb_4_l_fx_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15429\,
            lcout => if_generate_plus_mult1_un75_sum_axb_4_l_fx,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_rowlto2_sbtinv_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15297\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => un5_rowlto2_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \column_1_if_generate_plus_mult1_un75_sum_i_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15163\,
            lcout => \column_1_if_generate_plus_mult1_un75_sum_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16207\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15109\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15102\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHG_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16081\,
            in2 => \_gnd_net_\,
            in3 => \N__16414\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNIAGHGZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_4,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6Q_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16216\,
            in2 => \N__16411\,
            in3 => \N__16261\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNICK6QZ0\,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_5,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNITTA02_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__16235\,
            in1 => \N__16075\,
            in2 => \N__16060\,
            in3 => \N__16246\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un54_sum_axb_8,
            ltout => OPEN,
            carryin => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_6,
            carryout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EE_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16243\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIC9EEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQB_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16072\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI2FQBZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \un5_visiblex_cry_8_c_RNI1D62_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16210\,
            lcout => chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKN_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16073\,
            in2 => \_gnd_net_\,
            in3 => \N__16074\,
            lcout => \chessboardpixel_un152_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNI4UKNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
