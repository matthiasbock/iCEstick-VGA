// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 17 2015 19:42:52

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5947;
    wire N__5946;
    wire N__5945;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5929;
    wire N__5928;
    wire N__5927;
    wire N__5920;
    wire N__5919;
    wire N__5918;
    wire N__5911;
    wire N__5910;
    wire N__5909;
    wire N__5902;
    wire N__5901;
    wire N__5900;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5876;
    wire N__5875;
    wire N__5872;
    wire N__5871;
    wire N__5868;
    wire N__5867;
    wire N__5864;
    wire N__5855;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5832;
    wire N__5829;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5819;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5804;
    wire N__5799;
    wire N__5796;
    wire N__5793;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5781;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5769;
    wire N__5768;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5731;
    wire N__5730;
    wire N__5727;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5713;
    wire N__5710;
    wire N__5705;
    wire N__5704;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5683;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5655;
    wire N__5652;
    wire N__5649;
    wire N__5646;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5625;
    wire N__5624;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5601;
    wire N__5600;
    wire N__5599;
    wire N__5598;
    wire N__5597;
    wire N__5596;
    wire N__5595;
    wire N__5594;
    wire N__5593;
    wire N__5592;
    wire N__5591;
    wire N__5590;
    wire N__5589;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5540;
    wire N__5539;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5523;
    wire N__5522;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5485;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5459;
    wire N__5458;
    wire N__5457;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5449;
    wire N__5448;
    wire N__5447;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5400;
    wire N__5397;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5381;
    wire N__5378;
    wire N__5373;
    wire N__5368;
    wire N__5361;
    wire N__5352;
    wire N__5351;
    wire N__5350;
    wire N__5349;
    wire N__5348;
    wire N__5347;
    wire N__5346;
    wire N__5345;
    wire N__5340;
    wire N__5337;
    wire N__5330;
    wire N__5327;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5312;
    wire N__5309;
    wire N__5308;
    wire N__5307;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5293;
    wire N__5286;
    wire N__5277;
    wire N__5274;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5259;
    wire N__5256;
    wire N__5253;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5231;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5205;
    wire N__5200;
    wire N__5193;
    wire N__5190;
    wire N__5187;
    wire N__5184;
    wire N__5183;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5145;
    wire N__5144;
    wire N__5141;
    wire N__5140;
    wire N__5137;
    wire N__5136;
    wire N__5133;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5115;
    wire N__5112;
    wire N__5111;
    wire N__5108;
    wire N__5107;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5092;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5073;
    wire N__5070;
    wire N__5067;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5055;
    wire N__5054;
    wire N__5049;
    wire N__5046;
    wire N__5043;
    wire N__5040;
    wire N__5037;
    wire N__5034;
    wire N__5031;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5021;
    wire N__5020;
    wire N__5017;
    wire N__5016;
    wire N__5015;
    wire N__5012;
    wire N__5003;
    wire N__4998;
    wire N__4995;
    wire N__4992;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4977;
    wire N__4976;
    wire N__4973;
    wire N__4972;
    wire N__4971;
    wire N__4964;
    wire N__4961;
    wire N__4956;
    wire N__4953;
    wire N__4950;
    wire N__4947;
    wire N__4944;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4932;
    wire N__4929;
    wire N__4926;
    wire N__4925;
    wire N__4922;
    wire N__4921;
    wire N__4914;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4902;
    wire N__4899;
    wire N__4896;
    wire N__4893;
    wire N__4890;
    wire N__4887;
    wire N__4884;
    wire N__4881;
    wire N__4878;
    wire N__4875;
    wire N__4872;
    wire N__4869;
    wire N__4866;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4854;
    wire N__4851;
    wire N__4848;
    wire N__4847;
    wire N__4846;
    wire N__4845;
    wire N__4842;
    wire N__4839;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4821;
    wire N__4818;
    wire N__4815;
    wire N__4812;
    wire N__4809;
    wire N__4806;
    wire N__4803;
    wire N__4800;
    wire N__4797;
    wire N__4794;
    wire N__4791;
    wire N__4788;
    wire N__4785;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4773;
    wire N__4770;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4749;
    wire N__4746;
    wire N__4745;
    wire N__4742;
    wire N__4737;
    wire N__4734;
    wire N__4733;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4707;
    wire N__4704;
    wire N__4701;
    wire N__4698;
    wire N__4697;
    wire N__4694;
    wire N__4691;
    wire N__4686;
    wire N__4683;
    wire N__4680;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4665;
    wire N__4664;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4641;
    wire N__4640;
    wire N__4639;
    wire N__4636;
    wire N__4633;
    wire N__4632;
    wire N__4629;
    wire N__4620;
    wire N__4617;
    wire N__4614;
    wire N__4611;
    wire N__4610;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4593;
    wire N__4590;
    wire N__4587;
    wire N__4584;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4572;
    wire N__4571;
    wire N__4566;
    wire N__4563;
    wire N__4560;
    wire N__4559;
    wire N__4558;
    wire N__4557;
    wire N__4556;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4542;
    wire N__4539;
    wire N__4534;
    wire N__4533;
    wire N__4532;
    wire N__4527;
    wire N__4524;
    wire N__4519;
    wire N__4512;
    wire N__4509;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4491;
    wire N__4490;
    wire N__4489;
    wire N__4484;
    wire N__4481;
    wire N__4476;
    wire N__4475;
    wire N__4472;
    wire N__4471;
    wire N__4470;
    wire N__4469;
    wire N__4468;
    wire N__4467;
    wire N__4464;
    wire N__4461;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4447;
    wire N__4446;
    wire N__4443;
    wire N__4440;
    wire N__4435;
    wire N__4432;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4403;
    wire N__4392;
    wire N__4391;
    wire N__4386;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4371;
    wire N__4368;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4358;
    wire N__4357;
    wire N__4356;
    wire N__4353;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4341;
    wire N__4340;
    wire N__4339;
    wire N__4338;
    wire N__4337;
    wire N__4334;
    wire N__4327;
    wire N__4320;
    wire N__4317;
    wire N__4308;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4300;
    wire N__4299;
    wire N__4298;
    wire N__4297;
    wire N__4294;
    wire N__4291;
    wire N__4284;
    wire N__4281;
    wire N__4272;
    wire N__4269;
    wire N__4266;
    wire N__4263;
    wire N__4262;
    wire N__4261;
    wire N__4258;
    wire N__4257;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4230;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4218;
    wire N__4215;
    wire N__4214;
    wire N__4209;
    wire N__4206;
    wire N__4205;
    wire N__4200;
    wire N__4197;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4181;
    wire N__4180;
    wire N__4177;
    wire N__4176;
    wire N__4173;
    wire N__4170;
    wire N__4169;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4137;
    wire N__4136;
    wire N__4135;
    wire N__4134;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4126;
    wire N__4125;
    wire N__4124;
    wire N__4123;
    wire N__4120;
    wire N__4115;
    wire N__4110;
    wire N__4103;
    wire N__4102;
    wire N__4099;
    wire N__4094;
    wire N__4089;
    wire N__4086;
    wire N__4077;
    wire N__4076;
    wire N__4073;
    wire N__4072;
    wire N__4069;
    wire N__4068;
    wire N__4067;
    wire N__4066;
    wire N__4065;
    wire N__4062;
    wire N__4059;
    wire N__4056;
    wire N__4053;
    wire N__4050;
    wire N__4045;
    wire N__4042;
    wire N__4037;
    wire N__4026;
    wire N__4023;
    wire N__4022;
    wire N__4021;
    wire N__4020;
    wire N__4017;
    wire N__4016;
    wire N__4015;
    wire N__4010;
    wire N__4007;
    wire N__4006;
    wire N__4005;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3990;
    wire N__3987;
    wire N__3982;
    wire N__3969;
    wire N__3966;
    wire N__3963;
    wire N__3962;
    wire N__3961;
    wire N__3958;
    wire N__3957;
    wire N__3954;
    wire N__3953;
    wire N__3952;
    wire N__3949;
    wire N__3948;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3924;
    wire N__3909;
    wire N__3906;
    wire N__3905;
    wire N__3904;
    wire N__3903;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3888;
    wire N__3887;
    wire N__3886;
    wire N__3883;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3864;
    wire N__3861;
    wire N__3854;
    wire N__3843;
    wire N__3840;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3822;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3814;
    wire N__3813;
    wire N__3808;
    wire N__3805;
    wire N__3802;
    wire N__3799;
    wire N__3792;
    wire N__3789;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3777;
    wire N__3774;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3764;
    wire N__3763;
    wire N__3758;
    wire N__3755;
    wire N__3750;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3742;
    wire N__3737;
    wire N__3734;
    wire N__3729;
    wire N__3726;
    wire N__3723;
    wire N__3720;
    wire N__3717;
    wire N__3714;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3690;
    wire N__3689;
    wire N__3686;
    wire N__3685;
    wire N__3682;
    wire N__3681;
    wire N__3678;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3660;
    wire N__3657;
    wire N__3648;
    wire N__3645;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3633;
    wire N__3630;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3618;
    wire N__3615;
    wire N__3612;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3600;
    wire N__3597;
    wire N__3594;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3567;
    wire N__3566;
    wire N__3565;
    wire N__3562;
    wire N__3557;
    wire N__3552;
    wire N__3551;
    wire N__3546;
    wire N__3543;
    wire N__3540;
    wire N__3537;
    wire N__3536;
    wire N__3535;
    wire N__3528;
    wire N__3525;
    wire N__3522;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3509;
    wire N__3504;
    wire N__3503;
    wire N__3502;
    wire N__3501;
    wire N__3498;
    wire N__3495;
    wire N__3490;
    wire N__3483;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3471;
    wire N__3468;
    wire N__3465;
    wire N__3462;
    wire N__3459;
    wire N__3456;
    wire N__3453;
    wire N__3450;
    wire N__3447;
    wire N__3444;
    wire N__3441;
    wire N__3438;
    wire N__3435;
    wire N__3432;
    wire N__3429;
    wire N__3428;
    wire N__3427;
    wire N__3424;
    wire N__3421;
    wire N__3418;
    wire N__3411;
    wire N__3408;
    wire N__3405;
    wire N__3402;
    wire N__3399;
    wire N__3396;
    wire N__3393;
    wire N__3390;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3375;
    wire N__3372;
    wire N__3369;
    wire N__3366;
    wire N__3363;
    wire N__3360;
    wire N__3357;
    wire N__3356;
    wire N__3353;
    wire N__3350;
    wire N__3345;
    wire N__3342;
    wire N__3339;
    wire N__3336;
    wire N__3333;
    wire N__3330;
    wire N__3327;
    wire N__3324;
    wire N__3321;
    wire N__3318;
    wire N__3317;
    wire N__3316;
    wire N__3309;
    wire N__3306;
    wire N__3305;
    wire N__3304;
    wire N__3297;
    wire N__3294;
    wire N__3291;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3279;
    wire N__3276;
    wire N__3273;
    wire N__3272;
    wire N__3267;
    wire N__3264;
    wire N__3261;
    wire N__3258;
    wire N__3255;
    wire N__3252;
    wire N__3249;
    wire N__3246;
    wire N__3243;
    wire N__3240;
    wire N__3237;
    wire N__3234;
    wire N__3231;
    wire N__3228;
    wire N__3225;
    wire N__3222;
    wire N__3221;
    wire N__3216;
    wire N__3213;
    wire N__3212;
    wire N__3207;
    wire N__3204;
    wire N__3203;
    wire N__3200;
    wire N__3197;
    wire N__3192;
    wire N__3191;
    wire N__3190;
    wire N__3189;
    wire N__3188;
    wire N__3187;
    wire N__3186;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3166;
    wire N__3159;
    wire N__3158;
    wire N__3157;
    wire N__3156;
    wire N__3155;
    wire N__3154;
    wire N__3151;
    wire N__3144;
    wire N__3141;
    wire N__3138;
    wire N__3129;
    wire N__3126;
    wire N__3125;
    wire N__3124;
    wire N__3123;
    wire N__3120;
    wire N__3117;
    wire N__3114;
    wire N__3111;
    wire N__3102;
    wire N__3099;
    wire N__3098;
    wire N__3095;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3087;
    wire N__3084;
    wire N__3081;
    wire N__3078;
    wire N__3075;
    wire N__3066;
    wire N__3063;
    wire N__3060;
    wire N__3057;
    wire N__3054;
    wire N__3051;
    wire N__3048;
    wire N__3045;
    wire N__3042;
    wire N__3039;
    wire N__3036;
    wire N__3033;
    wire N__3030;
    wire N__3029;
    wire N__3028;
    wire N__3023;
    wire N__3022;
    wire N__3019;
    wire N__3016;
    wire N__3013;
    wire N__3010;
    wire N__3007;
    wire N__3000;
    wire N__2999;
    wire N__2998;
    wire N__2991;
    wire N__2988;
    wire N__2985;
    wire N__2982;
    wire N__2979;
    wire N__2976;
    wire N__2975;
    wire N__2974;
    wire N__2969;
    wire N__2968;
    wire N__2965;
    wire N__2962;
    wire N__2959;
    wire N__2952;
    wire N__2949;
    wire N__2948;
    wire N__2947;
    wire N__2946;
    wire N__2943;
    wire N__2942;
    wire N__2939;
    wire N__2934;
    wire N__2931;
    wire N__2928;
    wire N__2919;
    wire N__2916;
    wire N__2915;
    wire N__2912;
    wire N__2911;
    wire N__2908;
    wire N__2907;
    wire N__2906;
    wire N__2905;
    wire N__2902;
    wire N__2899;
    wire N__2892;
    wire N__2889;
    wire N__2880;
    wire N__2877;
    wire N__2876;
    wire N__2875;
    wire N__2874;
    wire N__2873;
    wire N__2872;
    wire N__2869;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2844;
    wire N__2841;
    wire N__2840;
    wire N__2839;
    wire N__2838;
    wire N__2835;
    wire N__2834;
    wire N__2833;
    wire N__2830;
    wire N__2825;
    wire N__2822;
    wire N__2819;
    wire N__2816;
    wire N__2805;
    wire N__2802;
    wire N__2799;
    wire N__2796;
    wire N__2793;
    wire N__2790;
    wire N__2787;
    wire N__2784;
    wire N__2781;
    wire N__2778;
    wire N__2775;
    wire N__2774;
    wire N__2771;
    wire N__2768;
    wire N__2765;
    wire N__2762;
    wire N__2759;
    wire N__2756;
    wire N__2753;
    wire N__2750;
    wire N__2745;
    wire N__2742;
    wire N__2739;
    wire N__2736;
    wire N__2733;
    wire N__2730;
    wire N__2727;
    wire N__2724;
    wire N__2721;
    wire N__2718;
    wire N__2715;
    wire N__2712;
    wire N__2709;
    wire N__2706;
    wire N__2703;
    wire N__2700;
    wire N__2697;
    wire N__2694;
    wire N__2691;
    wire N__2688;
    wire N__2685;
    wire N__2682;
    wire N__2679;
    wire N__2676;
    wire N__2673;
    wire N__2670;
    wire N__2667;
    wire N__2664;
    wire N__2661;
    wire N__2660;
    wire N__2655;
    wire N__2652;
    wire N__2649;
    wire N__2646;
    wire N__2643;
    wire N__2640;
    wire N__2637;
    wire N__2634;
    wire N__2631;
    wire N__2628;
    wire N__2625;
    wire \Clock50MHz.PixelClock ;
    wire Clock12MHz_c;
    wire VCCG0;
    wire GNDG0;
    wire un18_beamylto9_2_cascade_;
    wire un18_beamylt4;
    wire bfn_5_7_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire bfn_5_8_0_;
    wire un8_beamx_cry_9;
    wire bfn_6_2_0_;
    wire un20_beamy_cry_1;
    wire un20_beamy_cry_2;
    wire un20_beamy_cry_3;
    wire un20_beamy_cry_4;
    wire un20_beamy_cry_5;
    wire un20_beamy_cry_6;
    wire un20_beamy_cry_7;
    wire un20_beamy_cry_8;
    wire bfn_6_3_0_;
    wire un5_beamx_4_cascade_;
    wire beamY_RNI9DLCZ0Z_5_cascade_;
    wire un5_beamx_3;
    wire un5_beamx_2;
    wire un5_beamx_2_cascade_;
    wire un8_beamylto9_1_cascade_;
    wire un4_beamylt6_cascade_;
    wire un4_beamylt8_0_cascade_;
    wire un3_beamx_5;
    wire un3_beamx_7_cascade_;
    wire un1_beamxlt10_0_cascade_;
    wire HSync_c;
    wire un18_beamylt10_0;
    wire un8_beamy;
    wire un4_beamy_0;
    wire beamXZ0Z_10;
    wire un1_beamx_2;
    wire un13_beamylt7;
    wire un15_beamy_2_cascade_;
    wire bfn_6_7_0_;
    wire un5_visiblex_1_cry_0;
    wire beamXZ0Z_2;
    wire un5_visiblex_1_cry_1;
    wire beamXZ0Z_3;
    wire un5_visiblex_1_cry_2;
    wire beamXZ0Z_4;
    wire un5_visiblex_1_cry_3;
    wire beamXZ0Z_5;
    wire un5_visiblex_1_cry_4;
    wire beamXZ0Z_6;
    wire un5_visiblex_1_cry_5;
    wire beamXZ0Z_7;
    wire un5_visiblex_1_cry_6;
    wire un5_visiblex_1_cry_7;
    wire beamXZ0Z_8;
    wire bfn_6_8_0_;
    wire beamXZ0Z_9;
    wire un5_visiblex_1_cry_8;
    wire un5_visiblex_1_n_23_cascade_;
    wire bfn_7_2_0_;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_;
    wire beamY_fast_RNIGR79Z0Z_7_cascade_;
    wire beamY_RNIALEQ_0Z0Z_9;
    wire un20_beamy_cry_2_c_RNIBADZ0Z4;
    wire un20_beamy_cry_3_c_RNIDDEZ0Z4;
    wire un20_beamy_cry_6_c_RNIJMHZ0Z4;
    wire beamY_RNI9DLCZ0Z_5;
    wire un20_beamy_cry_4_c_RNIFGFZ0Z4;
    wire un13_visiblex_2_0;
    wire un12_visiblexlt9_0;
    wire un13_visiblex_0;
    wire font_un7_pixellt9_0;
    wire font_un14_pixellt9_0_cascade_;
    wire un13_visiblex_5;
    wire Pixel_0_sqmuxa_2;
    wire un13_visiblex_5_cascade_;
    wire un5_visiblex_1_n_31;
    wire un5_visiblex_1_n_30;
    wire N_159;
    wire bfn_7_7_0_;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1_cascade_;
    wire un5_visiblex_1_n_i_24;
    wire un5_visiblex_1_n_24;
    wire bfn_7_8_0_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3RZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4RZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_;
    wire un1_visiblex_if_generate_plus_mult1_un47_sum_i_8;
    wire un5_visiblex_1_n_23;
    wire un5_visiblex_1_cry_8_c_RNIHASCZ0Z_0;
    wire bfn_8_1_0_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_;
    wire un5_visibley_c3_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0Z_0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0;
    wire beamY_fastZ0Z_7;
    wire beamY_fastZ0Z_5;
    wire un5_visibley_c6_0_0_0;
    wire un5_visibley_c6_0_0_0_cascade_;
    wire un5_visibley_c3;
    wire beamY_RNIBV5PZ0Z_8;
    wire un13_visiblex_2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cascade_;
    wire beamY_fastZ0Z_3;
    wire beamY_fastZ0Z_4;
    wire un5_visibley_ac0_11_0_1_cascade_;
    wire beamY_fast_RNIGR79Z0Z_7;
    wire beamY_RNIALEQZ0Z_9;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cascade_;
    wire font_un11_pixellto9_7_0_cascade_;
    wire un8_beamx_cry_1_c_RNITP5AZ0;
    wire beamYZ0Z_0;
    wire font_un26_pixel_0_cascade_;
    wire un5_visibley_ac0_11_0_1;
    wire un5_visibley_c7;
    wire Pixel_0_sqmuxa_4;
    wire font_un11_pixel_0_7;
    wire un5_visibley_c7_cascade_;
    wire Pixel_0_sqmuxa_7;
    wire Pixel_0_sqmuxa_6;
    wire un15_beamy;
    wire Pixel_0_sqmuxa_7_cascade_;
    wire un13_visiblex_4;
    wire beamYZ0Z_4;
    wire beamYZ0Z_8;
    wire beamYZ0Z_7;
    wire beamYZ0Z_3;
    wire un1_beamylto9_1;
    wire beamYZ0Z_5;
    wire un1_beamylto9_2_cascade_;
    wire beamYZ0Z_9;
    wire VSync_c;
    wire un5_visiblex_1_n_26;
    wire bfn_8_6_0_;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKVZ0;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUDZ0Z1;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63_cascade_;
    wire beamXZ0Z_0;
    wire beamXZ0Z_1;
    wire beamX_RNIBKAZ0Z_1;
    wire un5_visiblex_1_n_25;
    wire un1_visiblex_if_generate_plus_mult1_un54_sum_i;
    wire bfn_9_1_0_;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250QZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIHZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_axb_6;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un40_sum;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_i_0;
    wire beamY_fastZ0Z_6;
    wire un20_beamy_cry_5_c_RNIHJGZ0Z4;
    wire beamYZ0Z_6;
    wire un20_beamy_cry_1_c_RNI97CZ0Z4;
    wire beamY_fastZ0Z_2;
    wire beamX_RNI5457Z0Z_5;
    wire bfn_9_5_0_;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_i;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05JZ0Z52;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEOZ0Z2;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63;
    wire un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBVZ0Z5;
    wire bfn_11_1_0_;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFVZ0Z81;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un47_sum;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_i_0;
    wire bfn_11_2_0_;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJZ0Z22;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_7;
    wire bfn_11_3_0_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONFZ0Z4;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEVZ0Z4;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBFZ0Z5;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6;
    wire un1_beamY_if_generate_plus_mult1_un61_sum;
    wire un1_beamY_if_generate_plus_mult1_un61_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un54_sum;
    wire un1_beamY_if_generate_plus_mult1_un54_sum_i_0;
    wire un1_visiblex_24;
    wire un19lto10_1_1_cascade_;
    wire un5_visiblex_1_n_28;
    wire bfn_11_5_0_;
    wire Pixel_1_RNOZ0Z_13;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOSZ0Z04;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVAZ0;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNPZ0Z5;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i_8;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8;
    wire un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7;
    wire Pixel_1_RNOZ0Z_6;
    wire un5_visiblex_1_n_27;
    wire un1_visiblex_if_generate_plus_mult1_un68_sum_i;
    wire CONSTANT_ONE_NET;
    wire beamYZ0Z_2;
    wire bfn_12_3_0_;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_2;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQZ0Z6;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85BZ0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_4;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LBZ0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_5;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_axb_7;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6;
    wire G_6_i_a4_0_0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0_cascade_;
    wire un1_beamY_if_generate_plus_mult1_un68_sum;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_i_0;
    wire un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0;
    wire beamY_i_2;
    wire un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0;
    wire beamYZ0Z_1;
    wire Pixel_1_RNOZ0Z_10;
    wire N_8_cascade_;
    wire N_11;
    wire un19_0_1;
    wire d_N_3_mux;
    wire un20_0_1_cascade_;
    wire Pixel_5_N_3_mux;
    wire Pixel_c;
    wire PixelClock_g;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__2634),
            .RESETB(N__5457),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__5956),
            .DIN(N__5955),
            .DOUT(N__5954),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__5956),
            .PADOUT(N__5955),
            .PADIN(N__5954),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5625),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__5947),
            .DIN(N__5946),
            .DOUT(N__5945),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__5947),
            .PADOUT(N__5946),
            .PADIN(N__5945),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3839),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__5938),
            .DIN(N__5937),
            .DOUT(N__5936),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__5938),
            .PADOUT(N__5937),
            .PADIN(N__5936),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2774),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__5929),
            .DIN(N__5928),
            .DOUT(N__5927),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__5929),
            .PADOUT(N__5928),
            .PADIN(N__5927),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3843),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__5920),
            .DIN(N__5919),
            .DOUT(N__5918),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__5920),
            .PADOUT(N__5919),
            .PADIN(N__5918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__5911),
            .DIN(N__5910),
            .DOUT(N__5909),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__5911),
            .PADOUT(N__5910),
            .PADIN(N__5909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2781),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__5902),
            .DIN(N__5901),
            .DOUT(N__5900),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__5902),
            .PADOUT(N__5901),
            .PADIN(N__5900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5624),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1314 (
            .O(N__5883),
            .I(N__5880));
    LocalMux I__1313 (
            .O(N__5880),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LBZ0));
    CascadeMux I__1312 (
            .O(N__5877),
            .I(N__5872));
    CascadeMux I__1311 (
            .O(N__5876),
            .I(N__5868));
    InMux I__1310 (
            .O(N__5875),
            .I(N__5864));
    InMux I__1309 (
            .O(N__5872),
            .I(N__5855));
    InMux I__1308 (
            .O(N__5871),
            .I(N__5855));
    InMux I__1307 (
            .O(N__5868),
            .I(N__5855));
    InMux I__1306 (
            .O(N__5867),
            .I(N__5855));
    LocalMux I__1305 (
            .O(N__5864),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0));
    LocalMux I__1304 (
            .O(N__5855),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0));
    CascadeMux I__1303 (
            .O(N__5850),
            .I(N__5847));
    InMux I__1302 (
            .O(N__5847),
            .I(N__5844));
    LocalMux I__1301 (
            .O(N__5844),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__1300 (
            .O(N__5841),
            .I(N__5838));
    LocalMux I__1299 (
            .O(N__5838),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__1298 (
            .O(N__5835),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6));
    InMux I__1297 (
            .O(N__5832),
            .I(N__5829));
    LocalMux I__1296 (
            .O(N__5829),
            .I(G_6_i_a4_0_0));
    CascadeMux I__1295 (
            .O(N__5826),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0_cascade_));
    InMux I__1294 (
            .O(N__5823),
            .I(N__5820));
    LocalMux I__1293 (
            .O(N__5820),
            .I(N__5815));
    InMux I__1292 (
            .O(N__5819),
            .I(N__5812));
    InMux I__1291 (
            .O(N__5818),
            .I(N__5809));
    Span4Mux_s0_h I__1290 (
            .O(N__5815),
            .I(N__5804));
    LocalMux I__1289 (
            .O(N__5812),
            .I(N__5804));
    LocalMux I__1288 (
            .O(N__5809),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    Odrv4 I__1287 (
            .O(N__5804),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum));
    InMux I__1286 (
            .O(N__5799),
            .I(N__5796));
    LocalMux I__1285 (
            .O(N__5796),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__1284 (
            .O(N__5793),
            .I(N__5789));
    InMux I__1283 (
            .O(N__5792),
            .I(N__5786));
    LocalMux I__1282 (
            .O(N__5789),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0));
    LocalMux I__1281 (
            .O(N__5786),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0));
    InMux I__1280 (
            .O(N__5781),
            .I(N__5777));
    InMux I__1279 (
            .O(N__5780),
            .I(N__5774));
    LocalMux I__1278 (
            .O(N__5777),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0));
    LocalMux I__1277 (
            .O(N__5774),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0));
    CascadeMux I__1276 (
            .O(N__5769),
            .I(N__5764));
    InMux I__1275 (
            .O(N__5768),
            .I(N__5761));
    InMux I__1274 (
            .O(N__5767),
            .I(N__5758));
    InMux I__1273 (
            .O(N__5764),
            .I(N__5755));
    LocalMux I__1272 (
            .O(N__5761),
            .I(N__5752));
    LocalMux I__1271 (
            .O(N__5758),
            .I(beamY_i_2));
    LocalMux I__1270 (
            .O(N__5755),
            .I(beamY_i_2));
    Odrv4 I__1269 (
            .O(N__5752),
            .I(beamY_i_2));
    InMux I__1268 (
            .O(N__5745),
            .I(N__5742));
    LocalMux I__1267 (
            .O(N__5742),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0));
    InMux I__1266 (
            .O(N__5739),
            .I(N__5735));
    InMux I__1265 (
            .O(N__5738),
            .I(N__5732));
    LocalMux I__1264 (
            .O(N__5735),
            .I(N__5727));
    LocalMux I__1263 (
            .O(N__5732),
            .I(N__5723));
    InMux I__1262 (
            .O(N__5731),
            .I(N__5720));
    CascadeMux I__1261 (
            .O(N__5730),
            .I(N__5717));
    Span4Mux_s1_h I__1260 (
            .O(N__5727),
            .I(N__5714));
    InMux I__1259 (
            .O(N__5726),
            .I(N__5710));
    Span4Mux_s2_h I__1258 (
            .O(N__5723),
            .I(N__5705));
    LocalMux I__1257 (
            .O(N__5720),
            .I(N__5705));
    InMux I__1256 (
            .O(N__5717),
            .I(N__5700));
    Span4Mux_h I__1255 (
            .O(N__5714),
            .I(N__5697));
    InMux I__1254 (
            .O(N__5713),
            .I(N__5694));
    LocalMux I__1253 (
            .O(N__5710),
            .I(N__5691));
    Span4Mux_h I__1252 (
            .O(N__5705),
            .I(N__5688));
    InMux I__1251 (
            .O(N__5704),
            .I(N__5683));
    InMux I__1250 (
            .O(N__5703),
            .I(N__5683));
    LocalMux I__1249 (
            .O(N__5700),
            .I(beamYZ0Z_1));
    Odrv4 I__1248 (
            .O(N__5697),
            .I(beamYZ0Z_1));
    LocalMux I__1247 (
            .O(N__5694),
            .I(beamYZ0Z_1));
    Odrv12 I__1246 (
            .O(N__5691),
            .I(beamYZ0Z_1));
    Odrv4 I__1245 (
            .O(N__5688),
            .I(beamYZ0Z_1));
    LocalMux I__1244 (
            .O(N__5683),
            .I(beamYZ0Z_1));
    InMux I__1243 (
            .O(N__5670),
            .I(N__5667));
    LocalMux I__1242 (
            .O(N__5667),
            .I(Pixel_1_RNOZ0Z_10));
    CascadeMux I__1241 (
            .O(N__5664),
            .I(N_8_cascade_));
    InMux I__1240 (
            .O(N__5661),
            .I(N__5658));
    LocalMux I__1239 (
            .O(N__5658),
            .I(N_11));
    InMux I__1238 (
            .O(N__5655),
            .I(N__5652));
    LocalMux I__1237 (
            .O(N__5652),
            .I(un19_0_1));
    InMux I__1236 (
            .O(N__5649),
            .I(N__5646));
    LocalMux I__1235 (
            .O(N__5646),
            .I(N__5643));
    Span4Mux_s1_h I__1234 (
            .O(N__5643),
            .I(N__5640));
    Odrv4 I__1233 (
            .O(N__5640),
            .I(d_N_3_mux));
    CascadeMux I__1232 (
            .O(N__5637),
            .I(un20_0_1_cascade_));
    InMux I__1231 (
            .O(N__5634),
            .I(N__5631));
    LocalMux I__1230 (
            .O(N__5631),
            .I(N__5628));
    Odrv12 I__1229 (
            .O(N__5628),
            .I(Pixel_5_N_3_mux));
    IoInMux I__1228 (
            .O(N__5625),
            .I(N__5621));
    IoInMux I__1227 (
            .O(N__5624),
            .I(N__5618));
    LocalMux I__1226 (
            .O(N__5621),
            .I(N__5615));
    LocalMux I__1225 (
            .O(N__5618),
            .I(N__5612));
    Span12Mux_s2_v I__1224 (
            .O(N__5615),
            .I(N__5609));
    Span4Mux_s3_v I__1223 (
            .O(N__5612),
            .I(N__5606));
    Odrv12 I__1222 (
            .O(N__5609),
            .I(Pixel_c));
    Odrv4 I__1221 (
            .O(N__5606),
            .I(Pixel_c));
    ClkMux I__1220 (
            .O(N__5601),
            .I(N__5562));
    ClkMux I__1219 (
            .O(N__5600),
            .I(N__5562));
    ClkMux I__1218 (
            .O(N__5599),
            .I(N__5562));
    ClkMux I__1217 (
            .O(N__5598),
            .I(N__5562));
    ClkMux I__1216 (
            .O(N__5597),
            .I(N__5562));
    ClkMux I__1215 (
            .O(N__5596),
            .I(N__5562));
    ClkMux I__1214 (
            .O(N__5595),
            .I(N__5562));
    ClkMux I__1213 (
            .O(N__5594),
            .I(N__5562));
    ClkMux I__1212 (
            .O(N__5593),
            .I(N__5562));
    ClkMux I__1211 (
            .O(N__5592),
            .I(N__5562));
    ClkMux I__1210 (
            .O(N__5591),
            .I(N__5562));
    ClkMux I__1209 (
            .O(N__5590),
            .I(N__5562));
    ClkMux I__1208 (
            .O(N__5589),
            .I(N__5562));
    GlobalMux I__1207 (
            .O(N__5562),
            .I(N__5559));
    gio2CtrlBuf I__1206 (
            .O(N__5559),
            .I(PixelClock_g));
    CascadeMux I__1205 (
            .O(N__5556),
            .I(N__5553));
    InMux I__1204 (
            .O(N__5553),
            .I(N__5550));
    LocalMux I__1203 (
            .O(N__5550),
            .I(N__5547));
    Odrv4 I__1202 (
            .O(N__5547),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNPZ0Z5));
    CascadeMux I__1201 (
            .O(N__5544),
            .I(N__5541));
    InMux I__1200 (
            .O(N__5541),
            .I(N__5534));
    InMux I__1199 (
            .O(N__5540),
            .I(N__5534));
    InMux I__1198 (
            .O(N__5539),
            .I(N__5531));
    LocalMux I__1197 (
            .O(N__5534),
            .I(N__5528));
    LocalMux I__1196 (
            .O(N__5531),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6));
    Odrv4 I__1195 (
            .O(N__5528),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6));
    InMux I__1194 (
            .O(N__5523),
            .I(N__5517));
    InMux I__1193 (
            .O(N__5522),
            .I(N__5517));
    LocalMux I__1192 (
            .O(N__5517),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__1191 (
            .O(N__5514),
            .I(N__5511));
    LocalMux I__1190 (
            .O(N__5511),
            .I(N__5508));
    Odrv4 I__1189 (
            .O(N__5508),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__1188 (
            .O(N__5505),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7));
    InMux I__1187 (
            .O(N__5502),
            .I(N__5499));
    LocalMux I__1186 (
            .O(N__5499),
            .I(Pixel_1_RNOZ0Z_6));
    InMux I__1185 (
            .O(N__5496),
            .I(N__5493));
    LocalMux I__1184 (
            .O(N__5493),
            .I(N__5489));
    InMux I__1183 (
            .O(N__5492),
            .I(N__5486));
    Span4Mux_s2_h I__1182 (
            .O(N__5489),
            .I(N__5480));
    LocalMux I__1181 (
            .O(N__5486),
            .I(N__5480));
    InMux I__1180 (
            .O(N__5485),
            .I(N__5477));
    Span4Mux_h I__1179 (
            .O(N__5480),
            .I(N__5474));
    LocalMux I__1178 (
            .O(N__5477),
            .I(un5_visiblex_1_n_27));
    Odrv4 I__1177 (
            .O(N__5474),
            .I(un5_visiblex_1_n_27));
    CascadeMux I__1176 (
            .O(N__5469),
            .I(N__5466));
    InMux I__1175 (
            .O(N__5466),
            .I(N__5463));
    LocalMux I__1174 (
            .O(N__5463),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_i));
    CascadeMux I__1173 (
            .O(N__5460),
            .I(N__5453));
    CascadeMux I__1172 (
            .O(N__5459),
            .I(N__5450));
    CascadeMux I__1171 (
            .O(N__5458),
            .I(N__5444));
    IoInMux I__1170 (
            .O(N__5457),
            .I(N__5439));
    InMux I__1169 (
            .O(N__5456),
            .I(N__5436));
    InMux I__1168 (
            .O(N__5453),
            .I(N__5433));
    InMux I__1167 (
            .O(N__5450),
            .I(N__5430));
    CascadeMux I__1166 (
            .O(N__5449),
            .I(N__5427));
    CascadeMux I__1165 (
            .O(N__5448),
            .I(N__5424));
    CascadeMux I__1164 (
            .O(N__5447),
            .I(N__5421));
    InMux I__1163 (
            .O(N__5444),
            .I(N__5418));
    CascadeMux I__1162 (
            .O(N__5443),
            .I(N__5415));
    CascadeMux I__1161 (
            .O(N__5442),
            .I(N__5412));
    LocalMux I__1160 (
            .O(N__5439),
            .I(N__5408));
    LocalMux I__1159 (
            .O(N__5436),
            .I(N__5405));
    LocalMux I__1158 (
            .O(N__5433),
            .I(N__5400));
    LocalMux I__1157 (
            .O(N__5430),
            .I(N__5400));
    InMux I__1156 (
            .O(N__5427),
            .I(N__5397));
    InMux I__1155 (
            .O(N__5424),
            .I(N__5392));
    InMux I__1154 (
            .O(N__5421),
            .I(N__5392));
    LocalMux I__1153 (
            .O(N__5418),
            .I(N__5389));
    InMux I__1152 (
            .O(N__5415),
            .I(N__5386));
    InMux I__1151 (
            .O(N__5412),
            .I(N__5381));
    InMux I__1150 (
            .O(N__5411),
            .I(N__5381));
    Span12Mux_s3_v I__1149 (
            .O(N__5408),
            .I(N__5378));
    Span4Mux_v I__1148 (
            .O(N__5405),
            .I(N__5373));
    Span4Mux_v I__1147 (
            .O(N__5400),
            .I(N__5373));
    LocalMux I__1146 (
            .O(N__5397),
            .I(N__5368));
    LocalMux I__1145 (
            .O(N__5392),
            .I(N__5368));
    Sp12to4 I__1144 (
            .O(N__5389),
            .I(N__5361));
    LocalMux I__1143 (
            .O(N__5386),
            .I(N__5361));
    LocalMux I__1142 (
            .O(N__5381),
            .I(N__5361));
    Odrv12 I__1141 (
            .O(N__5378),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1140 (
            .O(N__5373),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1139 (
            .O(N__5368),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1138 (
            .O(N__5361),
            .I(CONSTANT_ONE_NET));
    InMux I__1137 (
            .O(N__5352),
            .I(N__5340));
    InMux I__1136 (
            .O(N__5351),
            .I(N__5340));
    InMux I__1135 (
            .O(N__5350),
            .I(N__5337));
    InMux I__1134 (
            .O(N__5349),
            .I(N__5330));
    InMux I__1133 (
            .O(N__5348),
            .I(N__5330));
    InMux I__1132 (
            .O(N__5347),
            .I(N__5330));
    InMux I__1131 (
            .O(N__5346),
            .I(N__5327));
    InMux I__1130 (
            .O(N__5345),
            .I(N__5323));
    LocalMux I__1129 (
            .O(N__5340),
            .I(N__5320));
    LocalMux I__1128 (
            .O(N__5337),
            .I(N__5317));
    LocalMux I__1127 (
            .O(N__5330),
            .I(N__5312));
    LocalMux I__1126 (
            .O(N__5327),
            .I(N__5312));
    InMux I__1125 (
            .O(N__5326),
            .I(N__5309));
    LocalMux I__1124 (
            .O(N__5323),
            .I(N__5303));
    Span4Mux_h I__1123 (
            .O(N__5320),
            .I(N__5300));
    Span4Mux_s3_h I__1122 (
            .O(N__5317),
            .I(N__5293));
    Span4Mux_h I__1121 (
            .O(N__5312),
            .I(N__5293));
    LocalMux I__1120 (
            .O(N__5309),
            .I(N__5293));
    InMux I__1119 (
            .O(N__5308),
            .I(N__5286));
    InMux I__1118 (
            .O(N__5307),
            .I(N__5286));
    InMux I__1117 (
            .O(N__5306),
            .I(N__5286));
    Odrv12 I__1116 (
            .O(N__5303),
            .I(beamYZ0Z_2));
    Odrv4 I__1115 (
            .O(N__5300),
            .I(beamYZ0Z_2));
    Odrv4 I__1114 (
            .O(N__5293),
            .I(beamYZ0Z_2));
    LocalMux I__1113 (
            .O(N__5286),
            .I(beamYZ0Z_2));
    InMux I__1112 (
            .O(N__5277),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2));
    CascadeMux I__1111 (
            .O(N__5274),
            .I(N__5271));
    InMux I__1110 (
            .O(N__5271),
            .I(N__5268));
    LocalMux I__1109 (
            .O(N__5268),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQZ0Z6));
    InMux I__1108 (
            .O(N__5265),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__1107 (
            .O(N__5262),
            .I(N__5259));
    LocalMux I__1106 (
            .O(N__5259),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85BZ0));
    InMux I__1105 (
            .O(N__5256),
            .I(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__1104 (
            .O(N__5253),
            .I(N__5250));
    InMux I__1103 (
            .O(N__5250),
            .I(N__5247));
    LocalMux I__1102 (
            .O(N__5247),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__1101 (
            .O(N__5244),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1100 (
            .O(N__5241),
            .I(N__5238));
    LocalMux I__1099 (
            .O(N__5238),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__1098 (
            .O(N__5235),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__1097 (
            .O(N__5232),
            .I(N__5227));
    InMux I__1096 (
            .O(N__5231),
            .I(N__5224));
    InMux I__1095 (
            .O(N__5230),
            .I(N__5221));
    LocalMux I__1094 (
            .O(N__5227),
            .I(N__5217));
    LocalMux I__1093 (
            .O(N__5224),
            .I(N__5214));
    LocalMux I__1092 (
            .O(N__5221),
            .I(N__5211));
    InMux I__1091 (
            .O(N__5220),
            .I(N__5208));
    Span4Mux_s3_h I__1090 (
            .O(N__5217),
            .I(N__5205));
    Span4Mux_h I__1089 (
            .O(N__5214),
            .I(N__5200));
    Span4Mux_s3_h I__1088 (
            .O(N__5211),
            .I(N__5200));
    LocalMux I__1087 (
            .O(N__5208),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1086 (
            .O(N__5205),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    Odrv4 I__1085 (
            .O(N__5200),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum));
    CascadeMux I__1084 (
            .O(N__5193),
            .I(N__5190));
    InMux I__1083 (
            .O(N__5190),
            .I(N__5187));
    LocalMux I__1082 (
            .O(N__5187),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_i_0));
    InMux I__1081 (
            .O(N__5184),
            .I(N__5179));
    InMux I__1080 (
            .O(N__5183),
            .I(N__5176));
    InMux I__1079 (
            .O(N__5182),
            .I(N__5173));
    LocalMux I__1078 (
            .O(N__5179),
            .I(N__5170));
    LocalMux I__1077 (
            .O(N__5176),
            .I(N__5167));
    LocalMux I__1076 (
            .O(N__5173),
            .I(N__5164));
    Span4Mux_s3_h I__1075 (
            .O(N__5170),
            .I(N__5161));
    Odrv4 I__1074 (
            .O(N__5167),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1073 (
            .O(N__5164),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    Odrv4 I__1072 (
            .O(N__5161),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum));
    CascadeMux I__1071 (
            .O(N__5154),
            .I(N__5151));
    InMux I__1070 (
            .O(N__5151),
            .I(N__5148));
    LocalMux I__1069 (
            .O(N__5148),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__1068 (
            .O(N__5145),
            .I(N__5141));
    CascadeMux I__1067 (
            .O(N__5144),
            .I(N__5137));
    LocalMux I__1066 (
            .O(N__5141),
            .I(N__5133));
    InMux I__1065 (
            .O(N__5140),
            .I(N__5126));
    InMux I__1064 (
            .O(N__5137),
            .I(N__5126));
    InMux I__1063 (
            .O(N__5136),
            .I(N__5126));
    Span12Mux_s6_v I__1062 (
            .O(N__5133),
            .I(N__5123));
    LocalMux I__1061 (
            .O(N__5126),
            .I(N__5120));
    Odrv12 I__1060 (
            .O(N__5123),
            .I(un1_visiblex_24));
    Odrv4 I__1059 (
            .O(N__5120),
            .I(un1_visiblex_24));
    CascadeMux I__1058 (
            .O(N__5115),
            .I(un19lto10_1_1_cascade_));
    CascadeMux I__1057 (
            .O(N__5112),
            .I(N__5108));
    InMux I__1056 (
            .O(N__5111),
            .I(N__5102));
    InMux I__1055 (
            .O(N__5108),
            .I(N__5102));
    InMux I__1054 (
            .O(N__5107),
            .I(N__5099));
    LocalMux I__1053 (
            .O(N__5102),
            .I(N__5096));
    LocalMux I__1052 (
            .O(N__5099),
            .I(N__5093));
    Span4Mux_v I__1051 (
            .O(N__5096),
            .I(N__5087));
    Span4Mux_s1_h I__1050 (
            .O(N__5093),
            .I(N__5087));
    CascadeMux I__1049 (
            .O(N__5092),
            .I(N__5084));
    Span4Mux_h I__1048 (
            .O(N__5087),
            .I(N__5081));
    InMux I__1047 (
            .O(N__5084),
            .I(N__5078));
    Odrv4 I__1046 (
            .O(N__5081),
            .I(un5_visiblex_1_n_28));
    LocalMux I__1045 (
            .O(N__5078),
            .I(un5_visiblex_1_n_28));
    InMux I__1044 (
            .O(N__5073),
            .I(N__5070));
    LocalMux I__1043 (
            .O(N__5070),
            .I(Pixel_1_RNOZ0Z_13));
    InMux I__1042 (
            .O(N__5067),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__1041 (
            .O(N__5064),
            .I(N__5061));
    LocalMux I__1040 (
            .O(N__5061),
            .I(N__5058));
    Odrv4 I__1039 (
            .O(N__5058),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOSZ0Z04));
    InMux I__1038 (
            .O(N__5055),
            .I(N__5049));
    InMux I__1037 (
            .O(N__5054),
            .I(N__5049));
    LocalMux I__1036 (
            .O(N__5049),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVAZ0));
    InMux I__1035 (
            .O(N__5046),
            .I(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__1034 (
            .O(N__5043),
            .I(N__5040));
    LocalMux I__1033 (
            .O(N__5040),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJZ0Z22));
    InMux I__1032 (
            .O(N__5037),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__1031 (
            .O(N__5034),
            .I(N__5031));
    LocalMux I__1030 (
            .O(N__5031),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__1029 (
            .O(N__5028),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__1028 (
            .O(N__5025),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6_cascade_));
    CascadeMux I__1027 (
            .O(N__5022),
            .I(N__5017));
    InMux I__1026 (
            .O(N__5021),
            .I(N__5012));
    InMux I__1025 (
            .O(N__5020),
            .I(N__5003));
    InMux I__1024 (
            .O(N__5017),
            .I(N__5003));
    InMux I__1023 (
            .O(N__5016),
            .I(N__5003));
    InMux I__1022 (
            .O(N__5015),
            .I(N__5003));
    LocalMux I__1021 (
            .O(N__5012),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3));
    LocalMux I__1020 (
            .O(N__5003),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3));
    CascadeMux I__1019 (
            .O(N__4998),
            .I(N__4995));
    InMux I__1018 (
            .O(N__4995),
            .I(N__4992));
    LocalMux I__1017 (
            .O(N__4992),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__1016 (
            .O(N__4989),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__1015 (
            .O(N__4986),
            .I(N__4983));
    LocalMux I__1014 (
            .O(N__4983),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONFZ0Z4));
    InMux I__1013 (
            .O(N__4980),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__1012 (
            .O(N__4977),
            .I(N__4973));
    InMux I__1011 (
            .O(N__4976),
            .I(N__4964));
    InMux I__1010 (
            .O(N__4973),
            .I(N__4964));
    InMux I__1009 (
            .O(N__4972),
            .I(N__4964));
    InMux I__1008 (
            .O(N__4971),
            .I(N__4961));
    LocalMux I__1007 (
            .O(N__4964),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6));
    LocalMux I__1006 (
            .O(N__4961),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6));
    CascadeMux I__1005 (
            .O(N__4956),
            .I(N__4953));
    InMux I__1004 (
            .O(N__4953),
            .I(N__4950));
    LocalMux I__1003 (
            .O(N__4950),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEVZ0Z4));
    InMux I__1002 (
            .O(N__4947),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__1001 (
            .O(N__4944),
            .I(N__4941));
    LocalMux I__1000 (
            .O(N__4941),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBFZ0Z5));
    InMux I__999 (
            .O(N__4938),
            .I(N__4935));
    LocalMux I__998 (
            .O(N__4935),
            .I(N__4932));
    Odrv4 I__997 (
            .O(N__4932),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0));
    InMux I__996 (
            .O(N__4929),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3));
    CascadeMux I__995 (
            .O(N__4926),
            .I(N__4922));
    InMux I__994 (
            .O(N__4925),
            .I(N__4914));
    InMux I__993 (
            .O(N__4922),
            .I(N__4914));
    InMux I__992 (
            .O(N__4921),
            .I(N__4914));
    LocalMux I__991 (
            .O(N__4914),
            .I(N__4910));
    InMux I__990 (
            .O(N__4913),
            .I(N__4907));
    Odrv4 I__989 (
            .O(N__4910),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    LocalMux I__988 (
            .O(N__4907),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0));
    CascadeMux I__987 (
            .O(N__4902),
            .I(N__4899));
    InMux I__986 (
            .O(N__4899),
            .I(N__4896));
    LocalMux I__985 (
            .O(N__4896),
            .I(N__4893));
    Odrv4 I__984 (
            .O(N__4893),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFVZ0Z81));
    InMux I__983 (
            .O(N__4890),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__982 (
            .O(N__4887),
            .I(N__4884));
    LocalMux I__981 (
            .O(N__4884),
            .I(N__4881));
    Odrv4 I__980 (
            .O(N__4881),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1));
    CascadeMux I__979 (
            .O(N__4878),
            .I(N__4875));
    InMux I__978 (
            .O(N__4875),
            .I(N__4872));
    LocalMux I__977 (
            .O(N__4872),
            .I(N__4869));
    Odrv4 I__976 (
            .O(N__4869),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_7));
    InMux I__975 (
            .O(N__4866),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__974 (
            .O(N__4863),
            .I(N__4860));
    LocalMux I__973 (
            .O(N__4860),
            .I(N__4857));
    Odrv4 I__972 (
            .O(N__4857),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__971 (
            .O(N__4854),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__970 (
            .O(N__4851),
            .I(N__4848));
    LocalMux I__969 (
            .O(N__4848),
            .I(N__4842));
    CascadeMux I__968 (
            .O(N__4847),
            .I(N__4839));
    InMux I__967 (
            .O(N__4846),
            .I(N__4834));
    InMux I__966 (
            .O(N__4845),
            .I(N__4834));
    Span4Mux_s1_v I__965 (
            .O(N__4842),
            .I(N__4831));
    InMux I__964 (
            .O(N__4839),
            .I(N__4828));
    LocalMux I__963 (
            .O(N__4834),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    Odrv4 I__962 (
            .O(N__4831),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    LocalMux I__961 (
            .O(N__4828),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum));
    CascadeMux I__960 (
            .O(N__4821),
            .I(N__4818));
    InMux I__959 (
            .O(N__4818),
            .I(N__4815));
    LocalMux I__958 (
            .O(N__4815),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__957 (
            .O(N__4812),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__956 (
            .O(N__4809),
            .I(N__4806));
    LocalMux I__955 (
            .O(N__4806),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0));
    InMux I__954 (
            .O(N__4803),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3));
    CascadeMux I__953 (
            .O(N__4800),
            .I(N__4797));
    InMux I__952 (
            .O(N__4797),
            .I(N__4794));
    LocalMux I__951 (
            .O(N__4794),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1));
    InMux I__950 (
            .O(N__4791),
            .I(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__949 (
            .O(N__4788),
            .I(N__4785));
    LocalMux I__948 (
            .O(N__4785),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8));
    CascadeMux I__947 (
            .O(N__4782),
            .I(N__4779));
    InMux I__946 (
            .O(N__4779),
            .I(N__4776));
    LocalMux I__945 (
            .O(N__4776),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_i));
    InMux I__944 (
            .O(N__4773),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__943 (
            .O(N__4770),
            .I(N__4767));
    InMux I__942 (
            .O(N__4767),
            .I(N__4764));
    LocalMux I__941 (
            .O(N__4764),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05JZ0Z52));
    InMux I__940 (
            .O(N__4761),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__939 (
            .O(N__4758),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__938 (
            .O(N__4755),
            .I(N__4752));
    LocalMux I__937 (
            .O(N__4752),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__936 (
            .O(N__4749),
            .I(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7));
    CascadeMux I__935 (
            .O(N__4746),
            .I(N__4742));
    InMux I__934 (
            .O(N__4745),
            .I(N__4737));
    InMux I__933 (
            .O(N__4742),
            .I(N__4737));
    LocalMux I__932 (
            .O(N__4737),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEOZ0Z2));
    InMux I__931 (
            .O(N__4734),
            .I(N__4729));
    InMux I__930 (
            .O(N__4733),
            .I(N__4726));
    InMux I__929 (
            .O(N__4732),
            .I(N__4723));
    LocalMux I__928 (
            .O(N__4729),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63));
    LocalMux I__927 (
            .O(N__4726),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63));
    LocalMux I__926 (
            .O(N__4723),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63));
    InMux I__925 (
            .O(N__4716),
            .I(N__4713));
    LocalMux I__924 (
            .O(N__4713),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBVZ0Z5));
    InMux I__923 (
            .O(N__4710),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__922 (
            .O(N__4707),
            .I(N__4704));
    LocalMux I__921 (
            .O(N__4704),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51));
    InMux I__920 (
            .O(N__4701),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__919 (
            .O(N__4698),
            .I(N__4694));
    InMux I__918 (
            .O(N__4697),
            .I(N__4691));
    LocalMux I__917 (
            .O(N__4694),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51));
    LocalMux I__916 (
            .O(N__4691),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51));
    CascadeMux I__915 (
            .O(N__4686),
            .I(N__4683));
    InMux I__914 (
            .O(N__4683),
            .I(N__4680));
    LocalMux I__913 (
            .O(N__4680),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIHZ0Z1));
    InMux I__912 (
            .O(N__4677),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__911 (
            .O(N__4674),
            .I(N__4671));
    LocalMux I__910 (
            .O(N__4671),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__909 (
            .O(N__4668),
            .I(N__4665));
    LocalMux I__908 (
            .O(N__4665),
            .I(N__4660));
    CascadeMux I__907 (
            .O(N__4664),
            .I(N__4657));
    InMux I__906 (
            .O(N__4663),
            .I(N__4654));
    Span4Mux_s1_v I__905 (
            .O(N__4660),
            .I(N__4651));
    InMux I__904 (
            .O(N__4657),
            .I(N__4648));
    LocalMux I__903 (
            .O(N__4654),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    Odrv4 I__902 (
            .O(N__4651),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__901 (
            .O(N__4648),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6));
    CascadeMux I__900 (
            .O(N__4641),
            .I(N__4636));
    CascadeMux I__899 (
            .O(N__4640),
            .I(N__4633));
    CascadeMux I__898 (
            .O(N__4639),
            .I(N__4629));
    InMux I__897 (
            .O(N__4636),
            .I(N__4620));
    InMux I__896 (
            .O(N__4633),
            .I(N__4620));
    InMux I__895 (
            .O(N__4632),
            .I(N__4620));
    InMux I__894 (
            .O(N__4629),
            .I(N__4620));
    LocalMux I__893 (
            .O(N__4620),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0));
    InMux I__892 (
            .O(N__4617),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6));
    CascadeMux I__891 (
            .O(N__4614),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_));
    InMux I__890 (
            .O(N__4611),
            .I(N__4606));
    InMux I__889 (
            .O(N__4610),
            .I(N__4603));
    InMux I__888 (
            .O(N__4609),
            .I(N__4600));
    LocalMux I__887 (
            .O(N__4606),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    LocalMux I__886 (
            .O(N__4603),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    LocalMux I__885 (
            .O(N__4600),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum));
    InMux I__884 (
            .O(N__4593),
            .I(N__4590));
    LocalMux I__883 (
            .O(N__4590),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_i_0));
    CascadeMux I__882 (
            .O(N__4587),
            .I(N__4584));
    InMux I__881 (
            .O(N__4584),
            .I(N__4580));
    InMux I__880 (
            .O(N__4583),
            .I(N__4577));
    LocalMux I__879 (
            .O(N__4580),
            .I(beamY_fastZ0Z_6));
    LocalMux I__878 (
            .O(N__4577),
            .I(beamY_fastZ0Z_6));
    InMux I__877 (
            .O(N__4572),
            .I(N__4566));
    InMux I__876 (
            .O(N__4571),
            .I(N__4566));
    LocalMux I__875 (
            .O(N__4566),
            .I(N__4563));
    Odrv4 I__874 (
            .O(N__4563),
            .I(un20_beamy_cry_5_c_RNIHJGZ0Z4));
    InMux I__873 (
            .O(N__4560),
            .I(N__4551));
    InMux I__872 (
            .O(N__4559),
            .I(N__4551));
    InMux I__871 (
            .O(N__4558),
            .I(N__4548));
    InMux I__870 (
            .O(N__4557),
            .I(N__4545));
    InMux I__869 (
            .O(N__4556),
            .I(N__4542));
    LocalMux I__868 (
            .O(N__4551),
            .I(N__4539));
    LocalMux I__867 (
            .O(N__4548),
            .I(N__4534));
    LocalMux I__866 (
            .O(N__4545),
            .I(N__4534));
    LocalMux I__865 (
            .O(N__4542),
            .I(N__4527));
    Span4Mux_v I__864 (
            .O(N__4539),
            .I(N__4527));
    Span4Mux_h I__863 (
            .O(N__4534),
            .I(N__4524));
    InMux I__862 (
            .O(N__4533),
            .I(N__4519));
    InMux I__861 (
            .O(N__4532),
            .I(N__4519));
    Odrv4 I__860 (
            .O(N__4527),
            .I(beamYZ0Z_6));
    Odrv4 I__859 (
            .O(N__4524),
            .I(beamYZ0Z_6));
    LocalMux I__858 (
            .O(N__4519),
            .I(beamYZ0Z_6));
    InMux I__857 (
            .O(N__4512),
            .I(N__4509));
    LocalMux I__856 (
            .O(N__4509),
            .I(N__4505));
    InMux I__855 (
            .O(N__4508),
            .I(N__4502));
    Span4Mux_h I__854 (
            .O(N__4505),
            .I(N__4499));
    LocalMux I__853 (
            .O(N__4502),
            .I(N__4496));
    Odrv4 I__852 (
            .O(N__4499),
            .I(un20_beamy_cry_1_c_RNI97CZ0Z4));
    Odrv12 I__851 (
            .O(N__4496),
            .I(un20_beamy_cry_1_c_RNI97CZ0Z4));
    InMux I__850 (
            .O(N__4491),
            .I(N__4484));
    InMux I__849 (
            .O(N__4490),
            .I(N__4484));
    InMux I__848 (
            .O(N__4489),
            .I(N__4481));
    LocalMux I__847 (
            .O(N__4484),
            .I(beamY_fastZ0Z_2));
    LocalMux I__846 (
            .O(N__4481),
            .I(beamY_fastZ0Z_2));
    InMux I__845 (
            .O(N__4476),
            .I(N__4472));
    CEMux I__844 (
            .O(N__4475),
            .I(N__4464));
    LocalMux I__843 (
            .O(N__4472),
            .I(N__4461));
    InMux I__842 (
            .O(N__4471),
            .I(N__4458));
    CEMux I__841 (
            .O(N__4470),
            .I(N__4454));
    CEMux I__840 (
            .O(N__4469),
            .I(N__4451));
    CEMux I__839 (
            .O(N__4468),
            .I(N__4448));
    CEMux I__838 (
            .O(N__4467),
            .I(N__4443));
    LocalMux I__837 (
            .O(N__4464),
            .I(N__4440));
    Span4Mux_h I__836 (
            .O(N__4461),
            .I(N__4435));
    LocalMux I__835 (
            .O(N__4458),
            .I(N__4435));
    InMux I__834 (
            .O(N__4457),
            .I(N__4432));
    LocalMux I__833 (
            .O(N__4454),
            .I(N__4427));
    LocalMux I__832 (
            .O(N__4451),
            .I(N__4427));
    LocalMux I__831 (
            .O(N__4448),
            .I(N__4424));
    InMux I__830 (
            .O(N__4447),
            .I(N__4421));
    InMux I__829 (
            .O(N__4446),
            .I(N__4418));
    LocalMux I__828 (
            .O(N__4443),
            .I(N__4415));
    Span4Mux_h I__827 (
            .O(N__4440),
            .I(N__4412));
    Span4Mux_v I__826 (
            .O(N__4435),
            .I(N__4403));
    LocalMux I__825 (
            .O(N__4432),
            .I(N__4403));
    Span4Mux_h I__824 (
            .O(N__4427),
            .I(N__4403));
    Span4Mux_s2_v I__823 (
            .O(N__4424),
            .I(N__4403));
    LocalMux I__822 (
            .O(N__4421),
            .I(beamX_RNI5457Z0Z_5));
    LocalMux I__821 (
            .O(N__4418),
            .I(beamX_RNI5457Z0Z_5));
    Odrv12 I__820 (
            .O(N__4415),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__819 (
            .O(N__4412),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__818 (
            .O(N__4403),
            .I(beamX_RNI5457Z0Z_5));
    InMux I__817 (
            .O(N__4392),
            .I(N__4386));
    InMux I__816 (
            .O(N__4391),
            .I(N__4386));
    LocalMux I__815 (
            .O(N__4386),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__814 (
            .O(N__4383),
            .I(N__4380));
    InMux I__813 (
            .O(N__4380),
            .I(N__4377));
    LocalMux I__812 (
            .O(N__4377),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUDZ0Z1));
    InMux I__811 (
            .O(N__4374),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__810 (
            .O(N__4371),
            .I(N__4368));
    LocalMux I__809 (
            .O(N__4368),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__808 (
            .O(N__4365),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7));
    CascadeMux I__807 (
            .O(N__4362),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63_cascade_));
    CascadeMux I__806 (
            .O(N__4359),
            .I(N__4353));
    InMux I__805 (
            .O(N__4358),
            .I(N__4349));
    InMux I__804 (
            .O(N__4357),
            .I(N__4346));
    InMux I__803 (
            .O(N__4356),
            .I(N__4341));
    InMux I__802 (
            .O(N__4353),
            .I(N__4341));
    InMux I__801 (
            .O(N__4352),
            .I(N__4334));
    LocalMux I__800 (
            .O(N__4349),
            .I(N__4327));
    LocalMux I__799 (
            .O(N__4346),
            .I(N__4327));
    LocalMux I__798 (
            .O(N__4341),
            .I(N__4327));
    InMux I__797 (
            .O(N__4340),
            .I(N__4320));
    InMux I__796 (
            .O(N__4339),
            .I(N__4320));
    InMux I__795 (
            .O(N__4338),
            .I(N__4320));
    InMux I__794 (
            .O(N__4337),
            .I(N__4317));
    LocalMux I__793 (
            .O(N__4334),
            .I(beamXZ0Z_0));
    Odrv12 I__792 (
            .O(N__4327),
            .I(beamXZ0Z_0));
    LocalMux I__791 (
            .O(N__4320),
            .I(beamXZ0Z_0));
    LocalMux I__790 (
            .O(N__4317),
            .I(beamXZ0Z_0));
    InMux I__789 (
            .O(N__4308),
            .I(N__4304));
    CascadeMux I__788 (
            .O(N__4307),
            .I(N__4301));
    LocalMux I__787 (
            .O(N__4304),
            .I(N__4294));
    InMux I__786 (
            .O(N__4301),
            .I(N__4291));
    InMux I__785 (
            .O(N__4300),
            .I(N__4284));
    InMux I__784 (
            .O(N__4299),
            .I(N__4284));
    InMux I__783 (
            .O(N__4298),
            .I(N__4284));
    InMux I__782 (
            .O(N__4297),
            .I(N__4281));
    Odrv4 I__781 (
            .O(N__4294),
            .I(beamXZ0Z_1));
    LocalMux I__780 (
            .O(N__4291),
            .I(beamXZ0Z_1));
    LocalMux I__779 (
            .O(N__4284),
            .I(beamXZ0Z_1));
    LocalMux I__778 (
            .O(N__4281),
            .I(beamXZ0Z_1));
    InMux I__777 (
            .O(N__4272),
            .I(N__4269));
    LocalMux I__776 (
            .O(N__4269),
            .I(N__4266));
    Odrv4 I__775 (
            .O(N__4266),
            .I(beamX_RNIBKAZ0Z_1));
    InMux I__774 (
            .O(N__4263),
            .I(N__4258));
    InMux I__773 (
            .O(N__4262),
            .I(N__4252));
    InMux I__772 (
            .O(N__4261),
            .I(N__4252));
    LocalMux I__771 (
            .O(N__4258),
            .I(N__4249));
    InMux I__770 (
            .O(N__4257),
            .I(N__4246));
    LocalMux I__769 (
            .O(N__4252),
            .I(un5_visiblex_1_n_25));
    Odrv4 I__768 (
            .O(N__4249),
            .I(un5_visiblex_1_n_25));
    LocalMux I__767 (
            .O(N__4246),
            .I(un5_visiblex_1_n_25));
    CascadeMux I__766 (
            .O(N__4239),
            .I(N__4236));
    InMux I__765 (
            .O(N__4236),
            .I(N__4233));
    LocalMux I__764 (
            .O(N__4233),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_i));
    InMux I__763 (
            .O(N__4230),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2));
    CascadeMux I__762 (
            .O(N__4227),
            .I(N__4224));
    InMux I__761 (
            .O(N__4224),
            .I(N__4221));
    LocalMux I__760 (
            .O(N__4221),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250QZ0));
    InMux I__759 (
            .O(N__4218),
            .I(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__758 (
            .O(N__4215),
            .I(N__4209));
    InMux I__757 (
            .O(N__4214),
            .I(N__4209));
    LocalMux I__756 (
            .O(N__4209),
            .I(Pixel_0_sqmuxa_6));
    InMux I__755 (
            .O(N__4206),
            .I(N__4200));
    InMux I__754 (
            .O(N__4205),
            .I(N__4200));
    LocalMux I__753 (
            .O(N__4200),
            .I(N__4197));
    Span4Mux_h I__752 (
            .O(N__4197),
            .I(N__4194));
    Odrv4 I__751 (
            .O(N__4194),
            .I(un15_beamy));
    CascadeMux I__750 (
            .O(N__4191),
            .I(Pixel_0_sqmuxa_7_cascade_));
    InMux I__749 (
            .O(N__4188),
            .I(N__4185));
    LocalMux I__748 (
            .O(N__4185),
            .I(un13_visiblex_4));
    CascadeMux I__747 (
            .O(N__4182),
            .I(N__4177));
    InMux I__746 (
            .O(N__4181),
            .I(N__4173));
    InMux I__745 (
            .O(N__4180),
            .I(N__4170));
    InMux I__744 (
            .O(N__4177),
            .I(N__4165));
    InMux I__743 (
            .O(N__4176),
            .I(N__4162));
    LocalMux I__742 (
            .O(N__4173),
            .I(N__4157));
    LocalMux I__741 (
            .O(N__4170),
            .I(N__4157));
    InMux I__740 (
            .O(N__4169),
            .I(N__4154));
    InMux I__739 (
            .O(N__4168),
            .I(N__4151));
    LocalMux I__738 (
            .O(N__4165),
            .I(N__4148));
    LocalMux I__737 (
            .O(N__4162),
            .I(beamYZ0Z_4));
    Odrv4 I__736 (
            .O(N__4157),
            .I(beamYZ0Z_4));
    LocalMux I__735 (
            .O(N__4154),
            .I(beamYZ0Z_4));
    LocalMux I__734 (
            .O(N__4151),
            .I(beamYZ0Z_4));
    Odrv4 I__733 (
            .O(N__4148),
            .I(beamYZ0Z_4));
    InMux I__732 (
            .O(N__4137),
            .I(N__4130));
    InMux I__731 (
            .O(N__4136),
            .I(N__4127));
    InMux I__730 (
            .O(N__4135),
            .I(N__4120));
    InMux I__729 (
            .O(N__4134),
            .I(N__4115));
    InMux I__728 (
            .O(N__4133),
            .I(N__4115));
    LocalMux I__727 (
            .O(N__4130),
            .I(N__4110));
    LocalMux I__726 (
            .O(N__4127),
            .I(N__4110));
    InMux I__725 (
            .O(N__4126),
            .I(N__4103));
    InMux I__724 (
            .O(N__4125),
            .I(N__4103));
    InMux I__723 (
            .O(N__4124),
            .I(N__4103));
    InMux I__722 (
            .O(N__4123),
            .I(N__4099));
    LocalMux I__721 (
            .O(N__4120),
            .I(N__4094));
    LocalMux I__720 (
            .O(N__4115),
            .I(N__4094));
    Span4Mux_v I__719 (
            .O(N__4110),
            .I(N__4089));
    LocalMux I__718 (
            .O(N__4103),
            .I(N__4089));
    InMux I__717 (
            .O(N__4102),
            .I(N__4086));
    LocalMux I__716 (
            .O(N__4099),
            .I(beamYZ0Z_8));
    Odrv4 I__715 (
            .O(N__4094),
            .I(beamYZ0Z_8));
    Odrv4 I__714 (
            .O(N__4089),
            .I(beamYZ0Z_8));
    LocalMux I__713 (
            .O(N__4086),
            .I(beamYZ0Z_8));
    InMux I__712 (
            .O(N__4077),
            .I(N__4073));
    InMux I__711 (
            .O(N__4076),
            .I(N__4069));
    LocalMux I__710 (
            .O(N__4073),
            .I(N__4062));
    InMux I__709 (
            .O(N__4072),
            .I(N__4059));
    LocalMux I__708 (
            .O(N__4069),
            .I(N__4056));
    InMux I__707 (
            .O(N__4068),
            .I(N__4053));
    InMux I__706 (
            .O(N__4067),
            .I(N__4050));
    InMux I__705 (
            .O(N__4066),
            .I(N__4045));
    InMux I__704 (
            .O(N__4065),
            .I(N__4045));
    Span4Mux_h I__703 (
            .O(N__4062),
            .I(N__4042));
    LocalMux I__702 (
            .O(N__4059),
            .I(N__4037));
    Span4Mux_s1_v I__701 (
            .O(N__4056),
            .I(N__4037));
    LocalMux I__700 (
            .O(N__4053),
            .I(beamYZ0Z_7));
    LocalMux I__699 (
            .O(N__4050),
            .I(beamYZ0Z_7));
    LocalMux I__698 (
            .O(N__4045),
            .I(beamYZ0Z_7));
    Odrv4 I__697 (
            .O(N__4042),
            .I(beamYZ0Z_7));
    Odrv4 I__696 (
            .O(N__4037),
            .I(beamYZ0Z_7));
    CascadeMux I__695 (
            .O(N__4026),
            .I(N__4023));
    InMux I__694 (
            .O(N__4023),
            .I(N__4017));
    InMux I__693 (
            .O(N__4022),
            .I(N__4010));
    InMux I__692 (
            .O(N__4021),
            .I(N__4010));
    InMux I__691 (
            .O(N__4020),
            .I(N__4007));
    LocalMux I__690 (
            .O(N__4017),
            .I(N__4001));
    InMux I__689 (
            .O(N__4016),
            .I(N__3998));
    InMux I__688 (
            .O(N__4015),
            .I(N__3995));
    LocalMux I__687 (
            .O(N__4010),
            .I(N__3990));
    LocalMux I__686 (
            .O(N__4007),
            .I(N__3990));
    InMux I__685 (
            .O(N__4006),
            .I(N__3987));
    InMux I__684 (
            .O(N__4005),
            .I(N__3982));
    InMux I__683 (
            .O(N__4004),
            .I(N__3982));
    Odrv4 I__682 (
            .O(N__4001),
            .I(beamYZ0Z_3));
    LocalMux I__681 (
            .O(N__3998),
            .I(beamYZ0Z_3));
    LocalMux I__680 (
            .O(N__3995),
            .I(beamYZ0Z_3));
    Odrv4 I__679 (
            .O(N__3990),
            .I(beamYZ0Z_3));
    LocalMux I__678 (
            .O(N__3987),
            .I(beamYZ0Z_3));
    LocalMux I__677 (
            .O(N__3982),
            .I(beamYZ0Z_3));
    InMux I__676 (
            .O(N__3969),
            .I(N__3966));
    LocalMux I__675 (
            .O(N__3966),
            .I(un1_beamylto9_1));
    InMux I__674 (
            .O(N__3963),
            .I(N__3958));
    CascadeMux I__673 (
            .O(N__3962),
            .I(N__3954));
    InMux I__672 (
            .O(N__3961),
            .I(N__3949));
    LocalMux I__671 (
            .O(N__3958),
            .I(N__3944));
    InMux I__670 (
            .O(N__3957),
            .I(N__3941));
    InMux I__669 (
            .O(N__3954),
            .I(N__3938));
    InMux I__668 (
            .O(N__3953),
            .I(N__3933));
    InMux I__667 (
            .O(N__3952),
            .I(N__3933));
    LocalMux I__666 (
            .O(N__3949),
            .I(N__3930));
    InMux I__665 (
            .O(N__3948),
            .I(N__3927));
    InMux I__664 (
            .O(N__3947),
            .I(N__3924));
    Odrv4 I__663 (
            .O(N__3944),
            .I(beamYZ0Z_5));
    LocalMux I__662 (
            .O(N__3941),
            .I(beamYZ0Z_5));
    LocalMux I__661 (
            .O(N__3938),
            .I(beamYZ0Z_5));
    LocalMux I__660 (
            .O(N__3933),
            .I(beamYZ0Z_5));
    Odrv4 I__659 (
            .O(N__3930),
            .I(beamYZ0Z_5));
    LocalMux I__658 (
            .O(N__3927),
            .I(beamYZ0Z_5));
    LocalMux I__657 (
            .O(N__3924),
            .I(beamYZ0Z_5));
    CascadeMux I__656 (
            .O(N__3909),
            .I(un1_beamylto9_2_cascade_));
    InMux I__655 (
            .O(N__3906),
            .I(N__3899));
    InMux I__654 (
            .O(N__3905),
            .I(N__3896));
    InMux I__653 (
            .O(N__3904),
            .I(N__3892));
    InMux I__652 (
            .O(N__3903),
            .I(N__3889));
    InMux I__651 (
            .O(N__3902),
            .I(N__3883));
    LocalMux I__650 (
            .O(N__3899),
            .I(N__3878));
    LocalMux I__649 (
            .O(N__3896),
            .I(N__3878));
    InMux I__648 (
            .O(N__3895),
            .I(N__3875));
    LocalMux I__647 (
            .O(N__3892),
            .I(N__3872));
    LocalMux I__646 (
            .O(N__3889),
            .I(N__3869));
    InMux I__645 (
            .O(N__3888),
            .I(N__3864));
    InMux I__644 (
            .O(N__3887),
            .I(N__3864));
    InMux I__643 (
            .O(N__3886),
            .I(N__3861));
    LocalMux I__642 (
            .O(N__3883),
            .I(N__3854));
    Span4Mux_v I__641 (
            .O(N__3878),
            .I(N__3854));
    LocalMux I__640 (
            .O(N__3875),
            .I(N__3854));
    Odrv4 I__639 (
            .O(N__3872),
            .I(beamYZ0Z_9));
    Odrv4 I__638 (
            .O(N__3869),
            .I(beamYZ0Z_9));
    LocalMux I__637 (
            .O(N__3864),
            .I(beamYZ0Z_9));
    LocalMux I__636 (
            .O(N__3861),
            .I(beamYZ0Z_9));
    Odrv4 I__635 (
            .O(N__3854),
            .I(beamYZ0Z_9));
    IoInMux I__634 (
            .O(N__3843),
            .I(N__3840));
    LocalMux I__633 (
            .O(N__3840),
            .I(N__3836));
    IoInMux I__632 (
            .O(N__3839),
            .I(N__3833));
    Span12Mux_s11_v I__631 (
            .O(N__3836),
            .I(N__3830));
    LocalMux I__630 (
            .O(N__3833),
            .I(N__3827));
    Odrv12 I__629 (
            .O(N__3830),
            .I(VSync_c));
    Odrv12 I__628 (
            .O(N__3827),
            .I(VSync_c));
    InMux I__627 (
            .O(N__3822),
            .I(N__3818));
    InMux I__626 (
            .O(N__3821),
            .I(N__3815));
    LocalMux I__625 (
            .O(N__3818),
            .I(N__3808));
    LocalMux I__624 (
            .O(N__3815),
            .I(N__3808));
    InMux I__623 (
            .O(N__3814),
            .I(N__3805));
    InMux I__622 (
            .O(N__3813),
            .I(N__3802));
    Span4Mux_v I__621 (
            .O(N__3808),
            .I(N__3799));
    LocalMux I__620 (
            .O(N__3805),
            .I(un5_visiblex_1_n_26));
    LocalMux I__619 (
            .O(N__3802),
            .I(un5_visiblex_1_n_26));
    Odrv4 I__618 (
            .O(N__3799),
            .I(un5_visiblex_1_n_26));
    InMux I__617 (
            .O(N__3792),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__616 (
            .O(N__3789),
            .I(N__3785));
    InMux I__615 (
            .O(N__3788),
            .I(N__3782));
    LocalMux I__614 (
            .O(N__3785),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1));
    LocalMux I__613 (
            .O(N__3782),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1));
    CascadeMux I__612 (
            .O(N__3777),
            .I(N__3774));
    InMux I__611 (
            .O(N__3774),
            .I(N__3771));
    LocalMux I__610 (
            .O(N__3771),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKVZ0));
    InMux I__609 (
            .O(N__3768),
            .I(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__608 (
            .O(N__3765),
            .I(N__3758));
    InMux I__607 (
            .O(N__3764),
            .I(N__3758));
    InMux I__606 (
            .O(N__3763),
            .I(N__3755));
    LocalMux I__605 (
            .O(N__3758),
            .I(beamY_fastZ0Z_3));
    LocalMux I__604 (
            .O(N__3755),
            .I(beamY_fastZ0Z_3));
    CascadeMux I__603 (
            .O(N__3750),
            .I(N__3746));
    CascadeMux I__602 (
            .O(N__3749),
            .I(N__3743));
    InMux I__601 (
            .O(N__3746),
            .I(N__3737));
    InMux I__600 (
            .O(N__3743),
            .I(N__3737));
    InMux I__599 (
            .O(N__3742),
            .I(N__3734));
    LocalMux I__598 (
            .O(N__3737),
            .I(beamY_fastZ0Z_4));
    LocalMux I__597 (
            .O(N__3734),
            .I(beamY_fastZ0Z_4));
    CascadeMux I__596 (
            .O(N__3729),
            .I(un5_visibley_ac0_11_0_1_cascade_));
    InMux I__595 (
            .O(N__3726),
            .I(N__3723));
    LocalMux I__594 (
            .O(N__3723),
            .I(beamY_fast_RNIGR79Z0Z_7));
    InMux I__593 (
            .O(N__3720),
            .I(N__3717));
    LocalMux I__592 (
            .O(N__3717),
            .I(beamY_RNIALEQZ0Z_9));
    CascadeMux I__591 (
            .O(N__3714),
            .I(un1_beamY_if_generate_plus_mult1_un68_sum_cascade_));
    CascadeMux I__590 (
            .O(N__3711),
            .I(font_un11_pixellto9_7_0_cascade_));
    InMux I__589 (
            .O(N__3708),
            .I(N__3705));
    LocalMux I__588 (
            .O(N__3705),
            .I(N__3701));
    InMux I__587 (
            .O(N__3704),
            .I(N__3698));
    Span4Mux_h I__586 (
            .O(N__3701),
            .I(N__3695));
    LocalMux I__585 (
            .O(N__3698),
            .I(un8_beamx_cry_1_c_RNITP5AZ0));
    Odrv4 I__584 (
            .O(N__3695),
            .I(un8_beamx_cry_1_c_RNITP5AZ0));
    CascadeMux I__583 (
            .O(N__3690),
            .I(N__3686));
    CascadeMux I__582 (
            .O(N__3689),
            .I(N__3682));
    InMux I__581 (
            .O(N__3686),
            .I(N__3678));
    CascadeMux I__580 (
            .O(N__3685),
            .I(N__3674));
    InMux I__579 (
            .O(N__3682),
            .I(N__3671));
    InMux I__578 (
            .O(N__3681),
            .I(N__3668));
    LocalMux I__577 (
            .O(N__3678),
            .I(N__3665));
    InMux I__576 (
            .O(N__3677),
            .I(N__3660));
    InMux I__575 (
            .O(N__3674),
            .I(N__3660));
    LocalMux I__574 (
            .O(N__3671),
            .I(N__3657));
    LocalMux I__573 (
            .O(N__3668),
            .I(beamYZ0Z_0));
    Odrv4 I__572 (
            .O(N__3665),
            .I(beamYZ0Z_0));
    LocalMux I__571 (
            .O(N__3660),
            .I(beamYZ0Z_0));
    Odrv4 I__570 (
            .O(N__3657),
            .I(beamYZ0Z_0));
    CascadeMux I__569 (
            .O(N__3648),
            .I(font_un26_pixel_0_cascade_));
    InMux I__568 (
            .O(N__3645),
            .I(N__3641));
    InMux I__567 (
            .O(N__3644),
            .I(N__3638));
    LocalMux I__566 (
            .O(N__3641),
            .I(un5_visibley_ac0_11_0_1));
    LocalMux I__565 (
            .O(N__3638),
            .I(un5_visibley_ac0_11_0_1));
    CascadeMux I__564 (
            .O(N__3633),
            .I(N__3630));
    InMux I__563 (
            .O(N__3630),
            .I(N__3627));
    LocalMux I__562 (
            .O(N__3627),
            .I(un5_visibley_c7));
    InMux I__561 (
            .O(N__3624),
            .I(N__3621));
    LocalMux I__560 (
            .O(N__3621),
            .I(N__3618));
    Odrv4 I__559 (
            .O(N__3618),
            .I(Pixel_0_sqmuxa_4));
    InMux I__558 (
            .O(N__3615),
            .I(N__3612));
    LocalMux I__557 (
            .O(N__3612),
            .I(font_un11_pixel_0_7));
    CascadeMux I__556 (
            .O(N__3609),
            .I(un5_visibley_c7_cascade_));
    InMux I__555 (
            .O(N__3606),
            .I(N__3603));
    LocalMux I__554 (
            .O(N__3603),
            .I(Pixel_0_sqmuxa_7));
    CascadeMux I__553 (
            .O(N__3600),
            .I(un5_visibley_c3_cascade_));
    CascadeMux I__552 (
            .O(N__3597),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0Z_0_cascade_));
    CascadeMux I__551 (
            .O(N__3594),
            .I(N__3591));
    InMux I__550 (
            .O(N__3591),
            .I(N__3588));
    LocalMux I__549 (
            .O(N__3588),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0));
    CascadeMux I__548 (
            .O(N__3585),
            .I(N__3581));
    CascadeMux I__547 (
            .O(N__3584),
            .I(N__3578));
    InMux I__546 (
            .O(N__3581),
            .I(N__3575));
    InMux I__545 (
            .O(N__3578),
            .I(N__3572));
    LocalMux I__544 (
            .O(N__3575),
            .I(beamY_fastZ0Z_7));
    LocalMux I__543 (
            .O(N__3572),
            .I(beamY_fastZ0Z_7));
    InMux I__542 (
            .O(N__3567),
            .I(N__3562));
    InMux I__541 (
            .O(N__3566),
            .I(N__3557));
    InMux I__540 (
            .O(N__3565),
            .I(N__3557));
    LocalMux I__539 (
            .O(N__3562),
            .I(beamY_fastZ0Z_5));
    LocalMux I__538 (
            .O(N__3557),
            .I(beamY_fastZ0Z_5));
    InMux I__537 (
            .O(N__3552),
            .I(N__3546));
    InMux I__536 (
            .O(N__3551),
            .I(N__3546));
    LocalMux I__535 (
            .O(N__3546),
            .I(un5_visibley_c6_0_0_0));
    CascadeMux I__534 (
            .O(N__3543),
            .I(un5_visibley_c6_0_0_0_cascade_));
    CascadeMux I__533 (
            .O(N__3540),
            .I(N__3537));
    InMux I__532 (
            .O(N__3537),
            .I(N__3528));
    InMux I__531 (
            .O(N__3536),
            .I(N__3528));
    InMux I__530 (
            .O(N__3535),
            .I(N__3528));
    LocalMux I__529 (
            .O(N__3528),
            .I(un5_visibley_c3));
    InMux I__528 (
            .O(N__3525),
            .I(N__3522));
    LocalMux I__527 (
            .O(N__3522),
            .I(beamY_RNIBV5PZ0Z_8));
    InMux I__526 (
            .O(N__3519),
            .I(N__3516));
    LocalMux I__525 (
            .O(N__3516),
            .I(un13_visiblex_2));
    CascadeMux I__524 (
            .O(N__3513),
            .I(un1_beamY_if_generate_plus_mult1_un54_sum_cascade_));
    InMux I__523 (
            .O(N__3510),
            .I(N__3504));
    InMux I__522 (
            .O(N__3509),
            .I(N__3504));
    LocalMux I__521 (
            .O(N__3504),
            .I(N__3498));
    InMux I__520 (
            .O(N__3503),
            .I(N__3495));
    InMux I__519 (
            .O(N__3502),
            .I(N__3490));
    InMux I__518 (
            .O(N__3501),
            .I(N__3490));
    Odrv4 I__517 (
            .O(N__3498),
            .I(un5_visiblex_1_n_23));
    LocalMux I__516 (
            .O(N__3495),
            .I(un5_visiblex_1_n_23));
    LocalMux I__515 (
            .O(N__3490),
            .I(un5_visiblex_1_n_23));
    InMux I__514 (
            .O(N__3483),
            .I(N__3480));
    LocalMux I__513 (
            .O(N__3480),
            .I(un5_visiblex_1_cry_8_c_RNIHASCZ0Z_0));
    InMux I__512 (
            .O(N__3477),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2));
    InMux I__511 (
            .O(N__3474),
            .I(N__3471));
    LocalMux I__510 (
            .O(N__3471),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151));
    InMux I__509 (
            .O(N__3468),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__508 (
            .O(N__3465),
            .I(N__3462));
    LocalMux I__507 (
            .O(N__3462),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251));
    InMux I__506 (
            .O(N__3459),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__505 (
            .O(N__3456),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__504 (
            .O(N__3453),
            .I(N__3450));
    LocalMux I__503 (
            .O(N__3450),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    InMux I__502 (
            .O(N__3447),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__501 (
            .O(N__3444),
            .I(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_));
    CascadeMux I__500 (
            .O(N__3441),
            .I(N__3438));
    InMux I__499 (
            .O(N__3438),
            .I(N__3435));
    LocalMux I__498 (
            .O(N__3435),
            .I(un5_visiblex_1_n_i_24));
    InMux I__497 (
            .O(N__3432),
            .I(N__3429));
    LocalMux I__496 (
            .O(N__3429),
            .I(N__3424));
    InMux I__495 (
            .O(N__3428),
            .I(N__3421));
    InMux I__494 (
            .O(N__3427),
            .I(N__3418));
    Odrv4 I__493 (
            .O(N__3424),
            .I(un5_visiblex_1_n_24));
    LocalMux I__492 (
            .O(N__3421),
            .I(un5_visiblex_1_n_24));
    LocalMux I__491 (
            .O(N__3418),
            .I(un5_visiblex_1_n_24));
    InMux I__490 (
            .O(N__3411),
            .I(N__3408));
    LocalMux I__489 (
            .O(N__3408),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf));
    CascadeMux I__488 (
            .O(N__3405),
            .I(N__3402));
    InMux I__487 (
            .O(N__3402),
            .I(N__3399));
    LocalMux I__486 (
            .O(N__3399),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3RZ0));
    InMux I__485 (
            .O(N__3396),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__484 (
            .O(N__3393),
            .I(N__3390));
    InMux I__483 (
            .O(N__3390),
            .I(N__3387));
    LocalMux I__482 (
            .O(N__3387),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4RZ0));
    InMux I__481 (
            .O(N__3384),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5));
    CascadeMux I__480 (
            .O(N__3381),
            .I(N__3378));
    InMux I__479 (
            .O(N__3378),
            .I(N__3375));
    LocalMux I__478 (
            .O(N__3375),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO));
    InMux I__477 (
            .O(N__3372),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__476 (
            .O(N__3369),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__475 (
            .O(N__3366),
            .I(N__3363));
    LocalMux I__474 (
            .O(N__3363),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO));
    CascadeMux I__473 (
            .O(N__3360),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_));
    InMux I__472 (
            .O(N__3357),
            .I(N__3353));
    InMux I__471 (
            .O(N__3356),
            .I(N__3350));
    LocalMux I__470 (
            .O(N__3353),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0));
    LocalMux I__469 (
            .O(N__3350),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0));
    CascadeMux I__468 (
            .O(N__3345),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_));
    InMux I__467 (
            .O(N__3342),
            .I(N__3339));
    LocalMux I__466 (
            .O(N__3339),
            .I(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8));
    InMux I__465 (
            .O(N__3336),
            .I(N__3333));
    LocalMux I__464 (
            .O(N__3333),
            .I(un13_visiblex_5));
    InMux I__463 (
            .O(N__3330),
            .I(N__3327));
    LocalMux I__462 (
            .O(N__3327),
            .I(Pixel_0_sqmuxa_2));
    CascadeMux I__461 (
            .O(N__3324),
            .I(un13_visiblex_5_cascade_));
    CascadeMux I__460 (
            .O(N__3321),
            .I(N__3318));
    InMux I__459 (
            .O(N__3318),
            .I(N__3309));
    InMux I__458 (
            .O(N__3317),
            .I(N__3309));
    InMux I__457 (
            .O(N__3316),
            .I(N__3309));
    LocalMux I__456 (
            .O(N__3309),
            .I(un5_visiblex_1_n_31));
    InMux I__455 (
            .O(N__3306),
            .I(N__3297));
    InMux I__454 (
            .O(N__3305),
            .I(N__3297));
    InMux I__453 (
            .O(N__3304),
            .I(N__3297));
    LocalMux I__452 (
            .O(N__3297),
            .I(un5_visiblex_1_n_30));
    InMux I__451 (
            .O(N__3294),
            .I(N__3291));
    LocalMux I__450 (
            .O(N__3291),
            .I(N_159));
    InMux I__449 (
            .O(N__3288),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__448 (
            .O(N__3285),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__447 (
            .O(N__3282),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__446 (
            .O(N__3279),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7));
    CascadeMux I__445 (
            .O(N__3276),
            .I(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1_cascade_));
    InMux I__444 (
            .O(N__3273),
            .I(N__3267));
    InMux I__443 (
            .O(N__3272),
            .I(N__3267));
    LocalMux I__442 (
            .O(N__3267),
            .I(un20_beamy_cry_4_c_RNIFGFZ0Z4));
    InMux I__441 (
            .O(N__3264),
            .I(N__3261));
    LocalMux I__440 (
            .O(N__3261),
            .I(un13_visiblex_2_0));
    InMux I__439 (
            .O(N__3258),
            .I(N__3255));
    LocalMux I__438 (
            .O(N__3255),
            .I(un12_visiblexlt9_0));
    CascadeMux I__437 (
            .O(N__3252),
            .I(N__3249));
    InMux I__436 (
            .O(N__3249),
            .I(N__3246));
    LocalMux I__435 (
            .O(N__3246),
            .I(un13_visiblex_0));
    InMux I__434 (
            .O(N__3243),
            .I(N__3240));
    LocalMux I__433 (
            .O(N__3240),
            .I(font_un7_pixellt9_0));
    CascadeMux I__432 (
            .O(N__3237),
            .I(font_un14_pixellt9_0_cascade_));
    CascadeMux I__431 (
            .O(N__3234),
            .I(beamY_fast_RNIGR79Z0Z_7_cascade_));
    CascadeMux I__430 (
            .O(N__3231),
            .I(N__3228));
    InMux I__429 (
            .O(N__3228),
            .I(N__3225));
    LocalMux I__428 (
            .O(N__3225),
            .I(beamY_RNIALEQ_0Z0Z_9));
    InMux I__427 (
            .O(N__3222),
            .I(N__3216));
    InMux I__426 (
            .O(N__3221),
            .I(N__3216));
    LocalMux I__425 (
            .O(N__3216),
            .I(un20_beamy_cry_2_c_RNIBADZ0Z4));
    InMux I__424 (
            .O(N__3213),
            .I(N__3207));
    InMux I__423 (
            .O(N__3212),
            .I(N__3207));
    LocalMux I__422 (
            .O(N__3207),
            .I(un20_beamy_cry_3_c_RNIDDEZ0Z4));
    InMux I__421 (
            .O(N__3204),
            .I(N__3200));
    InMux I__420 (
            .O(N__3203),
            .I(N__3197));
    LocalMux I__419 (
            .O(N__3200),
            .I(un20_beamy_cry_6_c_RNIJMHZ0Z4));
    LocalMux I__418 (
            .O(N__3197),
            .I(un20_beamy_cry_6_c_RNIJMHZ0Z4));
    InMux I__417 (
            .O(N__3192),
            .I(N__3182));
    InMux I__416 (
            .O(N__3191),
            .I(N__3179));
    InMux I__415 (
            .O(N__3190),
            .I(N__3166));
    InMux I__414 (
            .O(N__3189),
            .I(N__3166));
    InMux I__413 (
            .O(N__3188),
            .I(N__3166));
    InMux I__412 (
            .O(N__3187),
            .I(N__3166));
    InMux I__411 (
            .O(N__3186),
            .I(N__3166));
    InMux I__410 (
            .O(N__3185),
            .I(N__3166));
    LocalMux I__409 (
            .O(N__3182),
            .I(beamY_RNI9DLCZ0Z_5));
    LocalMux I__408 (
            .O(N__3179),
            .I(beamY_RNI9DLCZ0Z_5));
    LocalMux I__407 (
            .O(N__3166),
            .I(beamY_RNI9DLCZ0Z_5));
    InMux I__406 (
            .O(N__3159),
            .I(N__3151));
    InMux I__405 (
            .O(N__3158),
            .I(N__3144));
    InMux I__404 (
            .O(N__3157),
            .I(N__3144));
    InMux I__403 (
            .O(N__3156),
            .I(N__3144));
    InMux I__402 (
            .O(N__3155),
            .I(N__3141));
    InMux I__401 (
            .O(N__3154),
            .I(N__3138));
    LocalMux I__400 (
            .O(N__3151),
            .I(beamXZ0Z_7));
    LocalMux I__399 (
            .O(N__3144),
            .I(beamXZ0Z_7));
    LocalMux I__398 (
            .O(N__3141),
            .I(beamXZ0Z_7));
    LocalMux I__397 (
            .O(N__3138),
            .I(beamXZ0Z_7));
    InMux I__396 (
            .O(N__3129),
            .I(un5_visiblex_1_cry_6));
    InMux I__395 (
            .O(N__3126),
            .I(N__3120));
    InMux I__394 (
            .O(N__3125),
            .I(N__3117));
    InMux I__393 (
            .O(N__3124),
            .I(N__3114));
    InMux I__392 (
            .O(N__3123),
            .I(N__3111));
    LocalMux I__391 (
            .O(N__3120),
            .I(beamXZ0Z_8));
    LocalMux I__390 (
            .O(N__3117),
            .I(beamXZ0Z_8));
    LocalMux I__389 (
            .O(N__3114),
            .I(beamXZ0Z_8));
    LocalMux I__388 (
            .O(N__3111),
            .I(beamXZ0Z_8));
    InMux I__387 (
            .O(N__3102),
            .I(bfn_6_8_0_));
    CascadeMux I__386 (
            .O(N__3099),
            .I(N__3095));
    InMux I__385 (
            .O(N__3098),
            .I(N__3091));
    InMux I__384 (
            .O(N__3095),
            .I(N__3088));
    InMux I__383 (
            .O(N__3094),
            .I(N__3084));
    LocalMux I__382 (
            .O(N__3091),
            .I(N__3081));
    LocalMux I__381 (
            .O(N__3088),
            .I(N__3078));
    InMux I__380 (
            .O(N__3087),
            .I(N__3075));
    LocalMux I__379 (
            .O(N__3084),
            .I(beamXZ0Z_9));
    Odrv4 I__378 (
            .O(N__3081),
            .I(beamXZ0Z_9));
    Odrv4 I__377 (
            .O(N__3078),
            .I(beamXZ0Z_9));
    LocalMux I__376 (
            .O(N__3075),
            .I(beamXZ0Z_9));
    InMux I__375 (
            .O(N__3066),
            .I(un5_visiblex_1_cry_8));
    CascadeMux I__374 (
            .O(N__3063),
            .I(un5_visiblex_1_n_23_cascade_));
    InMux I__373 (
            .O(N__3060),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__372 (
            .O(N__3057),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__371 (
            .O(N__3054),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5));
    CascadeMux I__370 (
            .O(N__3051),
            .I(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_));
    InMux I__369 (
            .O(N__3048),
            .I(N__3045));
    LocalMux I__368 (
            .O(N__3045),
            .I(N__3042));
    Odrv4 I__367 (
            .O(N__3042),
            .I(un8_beamy));
    CascadeMux I__366 (
            .O(N__3039),
            .I(N__3036));
    InMux I__365 (
            .O(N__3036),
            .I(N__3033));
    LocalMux I__364 (
            .O(N__3033),
            .I(un4_beamy_0));
    InMux I__363 (
            .O(N__3030),
            .I(N__3023));
    InMux I__362 (
            .O(N__3029),
            .I(N__3023));
    InMux I__361 (
            .O(N__3028),
            .I(N__3019));
    LocalMux I__360 (
            .O(N__3023),
            .I(N__3016));
    InMux I__359 (
            .O(N__3022),
            .I(N__3013));
    LocalMux I__358 (
            .O(N__3019),
            .I(N__3010));
    Span4Mux_h I__357 (
            .O(N__3016),
            .I(N__3007));
    LocalMux I__356 (
            .O(N__3013),
            .I(beamXZ0Z_10));
    Odrv4 I__355 (
            .O(N__3010),
            .I(beamXZ0Z_10));
    Odrv4 I__354 (
            .O(N__3007),
            .I(beamXZ0Z_10));
    InMux I__353 (
            .O(N__3000),
            .I(N__2991));
    InMux I__352 (
            .O(N__2999),
            .I(N__2991));
    InMux I__351 (
            .O(N__2998),
            .I(N__2991));
    LocalMux I__350 (
            .O(N__2991),
            .I(un1_beamx_2));
    InMux I__349 (
            .O(N__2988),
            .I(N__2985));
    LocalMux I__348 (
            .O(N__2985),
            .I(un13_beamylt7));
    CascadeMux I__347 (
            .O(N__2982),
            .I(un15_beamy_2_cascade_));
    InMux I__346 (
            .O(N__2979),
            .I(un5_visiblex_1_cry_0));
    InMux I__345 (
            .O(N__2976),
            .I(N__2969));
    InMux I__344 (
            .O(N__2975),
            .I(N__2969));
    InMux I__343 (
            .O(N__2974),
            .I(N__2965));
    LocalMux I__342 (
            .O(N__2969),
            .I(N__2962));
    InMux I__341 (
            .O(N__2968),
            .I(N__2959));
    LocalMux I__340 (
            .O(N__2965),
            .I(beamXZ0Z_2));
    Odrv4 I__339 (
            .O(N__2962),
            .I(beamXZ0Z_2));
    LocalMux I__338 (
            .O(N__2959),
            .I(beamXZ0Z_2));
    InMux I__337 (
            .O(N__2952),
            .I(un5_visiblex_1_cry_1));
    CascadeMux I__336 (
            .O(N__2949),
            .I(N__2943));
    InMux I__335 (
            .O(N__2948),
            .I(N__2939));
    InMux I__334 (
            .O(N__2947),
            .I(N__2934));
    InMux I__333 (
            .O(N__2946),
            .I(N__2934));
    InMux I__332 (
            .O(N__2943),
            .I(N__2931));
    InMux I__331 (
            .O(N__2942),
            .I(N__2928));
    LocalMux I__330 (
            .O(N__2939),
            .I(beamXZ0Z_3));
    LocalMux I__329 (
            .O(N__2934),
            .I(beamXZ0Z_3));
    LocalMux I__328 (
            .O(N__2931),
            .I(beamXZ0Z_3));
    LocalMux I__327 (
            .O(N__2928),
            .I(beamXZ0Z_3));
    InMux I__326 (
            .O(N__2919),
            .I(un5_visiblex_1_cry_2));
    CascadeMux I__325 (
            .O(N__2916),
            .I(N__2912));
    CascadeMux I__324 (
            .O(N__2915),
            .I(N__2908));
    InMux I__323 (
            .O(N__2912),
            .I(N__2902));
    InMux I__322 (
            .O(N__2911),
            .I(N__2899));
    InMux I__321 (
            .O(N__2908),
            .I(N__2892));
    InMux I__320 (
            .O(N__2907),
            .I(N__2892));
    InMux I__319 (
            .O(N__2906),
            .I(N__2892));
    InMux I__318 (
            .O(N__2905),
            .I(N__2889));
    LocalMux I__317 (
            .O(N__2902),
            .I(beamXZ0Z_4));
    LocalMux I__316 (
            .O(N__2899),
            .I(beamXZ0Z_4));
    LocalMux I__315 (
            .O(N__2892),
            .I(beamXZ0Z_4));
    LocalMux I__314 (
            .O(N__2889),
            .I(beamXZ0Z_4));
    InMux I__313 (
            .O(N__2880),
            .I(un5_visiblex_1_cry_3));
    InMux I__312 (
            .O(N__2877),
            .I(N__2869));
    InMux I__311 (
            .O(N__2876),
            .I(N__2864));
    InMux I__310 (
            .O(N__2875),
            .I(N__2864));
    InMux I__309 (
            .O(N__2874),
            .I(N__2861));
    InMux I__308 (
            .O(N__2873),
            .I(N__2858));
    InMux I__307 (
            .O(N__2872),
            .I(N__2855));
    LocalMux I__306 (
            .O(N__2869),
            .I(beamXZ0Z_5));
    LocalMux I__305 (
            .O(N__2864),
            .I(beamXZ0Z_5));
    LocalMux I__304 (
            .O(N__2861),
            .I(beamXZ0Z_5));
    LocalMux I__303 (
            .O(N__2858),
            .I(beamXZ0Z_5));
    LocalMux I__302 (
            .O(N__2855),
            .I(beamXZ0Z_5));
    InMux I__301 (
            .O(N__2844),
            .I(un5_visiblex_1_cry_4));
    CascadeMux I__300 (
            .O(N__2841),
            .I(N__2835));
    InMux I__299 (
            .O(N__2840),
            .I(N__2830));
    InMux I__298 (
            .O(N__2839),
            .I(N__2825));
    InMux I__297 (
            .O(N__2838),
            .I(N__2825));
    InMux I__296 (
            .O(N__2835),
            .I(N__2822));
    InMux I__295 (
            .O(N__2834),
            .I(N__2819));
    InMux I__294 (
            .O(N__2833),
            .I(N__2816));
    LocalMux I__293 (
            .O(N__2830),
            .I(beamXZ0Z_6));
    LocalMux I__292 (
            .O(N__2825),
            .I(beamXZ0Z_6));
    LocalMux I__291 (
            .O(N__2822),
            .I(beamXZ0Z_6));
    LocalMux I__290 (
            .O(N__2819),
            .I(beamXZ0Z_6));
    LocalMux I__289 (
            .O(N__2816),
            .I(beamXZ0Z_6));
    InMux I__288 (
            .O(N__2805),
            .I(un5_visiblex_1_cry_5));
    CascadeMux I__287 (
            .O(N__2802),
            .I(un4_beamylt6_cascade_));
    CascadeMux I__286 (
            .O(N__2799),
            .I(un4_beamylt8_0_cascade_));
    CascadeMux I__285 (
            .O(N__2796),
            .I(N__2793));
    InMux I__284 (
            .O(N__2793),
            .I(N__2790));
    LocalMux I__283 (
            .O(N__2790),
            .I(un3_beamx_5));
    CascadeMux I__282 (
            .O(N__2787),
            .I(un3_beamx_7_cascade_));
    CascadeMux I__281 (
            .O(N__2784),
            .I(un1_beamxlt10_0_cascade_));
    IoInMux I__280 (
            .O(N__2781),
            .I(N__2778));
    LocalMux I__279 (
            .O(N__2778),
            .I(N__2775));
    Span4Mux_s2_v I__278 (
            .O(N__2775),
            .I(N__2771));
    IoInMux I__277 (
            .O(N__2774),
            .I(N__2768));
    Span4Mux_h I__276 (
            .O(N__2771),
            .I(N__2765));
    LocalMux I__275 (
            .O(N__2768),
            .I(N__2762));
    Span4Mux_v I__274 (
            .O(N__2765),
            .I(N__2759));
    IoSpan4Mux I__273 (
            .O(N__2762),
            .I(N__2756));
    Span4Mux_v I__272 (
            .O(N__2759),
            .I(N__2753));
    Span4Mux_s3_v I__271 (
            .O(N__2756),
            .I(N__2750));
    Odrv4 I__270 (
            .O(N__2753),
            .I(HSync_c));
    Odrv4 I__269 (
            .O(N__2750),
            .I(HSync_c));
    InMux I__268 (
            .O(N__2745),
            .I(N__2742));
    LocalMux I__267 (
            .O(N__2742),
            .I(un18_beamylt10_0));
    InMux I__266 (
            .O(N__2739),
            .I(un20_beamy_cry_7));
    InMux I__265 (
            .O(N__2736),
            .I(bfn_6_3_0_));
    CascadeMux I__264 (
            .O(N__2733),
            .I(un5_beamx_4_cascade_));
    CascadeMux I__263 (
            .O(N__2730),
            .I(beamY_RNI9DLCZ0Z_5_cascade_));
    InMux I__262 (
            .O(N__2727),
            .I(N__2724));
    LocalMux I__261 (
            .O(N__2724),
            .I(un5_beamx_3));
    InMux I__260 (
            .O(N__2721),
            .I(N__2718));
    LocalMux I__259 (
            .O(N__2718),
            .I(un5_beamx_2));
    CascadeMux I__258 (
            .O(N__2715),
            .I(un5_beamx_2_cascade_));
    CascadeMux I__257 (
            .O(N__2712),
            .I(un8_beamylto9_1_cascade_));
    InMux I__256 (
            .O(N__2709),
            .I(un8_beamx_cry_9));
    InMux I__255 (
            .O(N__2706),
            .I(un20_beamy_cry_1));
    InMux I__254 (
            .O(N__2703),
            .I(un20_beamy_cry_2));
    InMux I__253 (
            .O(N__2700),
            .I(un20_beamy_cry_3));
    InMux I__252 (
            .O(N__2697),
            .I(un20_beamy_cry_4));
    InMux I__251 (
            .O(N__2694),
            .I(un20_beamy_cry_5));
    InMux I__250 (
            .O(N__2691),
            .I(un20_beamy_cry_6));
    InMux I__249 (
            .O(N__2688),
            .I(un8_beamx_cry_1));
    InMux I__248 (
            .O(N__2685),
            .I(un8_beamx_cry_2));
    InMux I__247 (
            .O(N__2682),
            .I(un8_beamx_cry_3));
    InMux I__246 (
            .O(N__2679),
            .I(un8_beamx_cry_4));
    InMux I__245 (
            .O(N__2676),
            .I(un8_beamx_cry_5));
    InMux I__244 (
            .O(N__2673),
            .I(un8_beamx_cry_6));
    InMux I__243 (
            .O(N__2670),
            .I(un8_beamx_cry_7));
    InMux I__242 (
            .O(N__2667),
            .I(bfn_5_8_0_));
    CascadeMux I__241 (
            .O(N__2664),
            .I(un18_beamylto9_2_cascade_));
    InMux I__240 (
            .O(N__2661),
            .I(N__2655));
    InMux I__239 (
            .O(N__2660),
            .I(N__2655));
    LocalMux I__238 (
            .O(N__2655),
            .I(un18_beamylt4));
    IoInMux I__237 (
            .O(N__2652),
            .I(N__2649));
    LocalMux I__236 (
            .O(N__2649),
            .I(N__2646));
    IoSpan4Mux I__235 (
            .O(N__2646),
            .I(N__2643));
    IoSpan4Mux I__234 (
            .O(N__2643),
            .I(N__2640));
    IoSpan4Mux I__233 (
            .O(N__2640),
            .I(N__2637));
    Odrv4 I__232 (
            .O(N__2637),
            .I(\Clock50MHz.PixelClock ));
    IoInMux I__231 (
            .O(N__2634),
            .I(N__2631));
    LocalMux I__230 (
            .O(N__2631),
            .I(N__2628));
    IoSpan4Mux I__229 (
            .O(N__2628),
            .I(N__2625));
    Odrv4 I__228 (
            .O(N__2625),
            .I(Clock12MHz_c));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(un5_visiblex_1_cry_7),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_6_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_2_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(un20_beamy_cry_8),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_1_0_));
    defparam IN_MUX_bfv_9_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_1_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_3_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__2652),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam beamX_RNIQCL_1_LC_5_6_0.C_ON=1'b0;
    defparam beamX_RNIQCL_1_LC_5_6_0.SEQ_MODE=4'b0000;
    defparam beamX_RNIQCL_1_LC_5_6_0.LUT_INIT=16'b0000011100001111;
    LogicCell40 beamX_RNIQCL_1_LC_5_6_0 (
            .in0(N__2975),
            .in1(N__4298),
            .in2(N__2949),
            .in3(N__4338),
            .lcout(un18_beamylt4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_5_6_1.C_ON=1'b0;
    defparam beamX_0_LC_5_6_1.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_5_6_1.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamX_0_LC_5_6_1 (
            .in0(N__4339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4447),
            .lcout(beamXZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5591),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_5_6_2.C_ON=1'b0;
    defparam beamX_1_LC_5_6_2.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_5_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 beamX_1_LC_5_6_2 (
            .in0(_gnd_net_),
            .in1(N__4300),
            .in2(_gnd_net_),
            .in3(N__4340),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5591),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNII5M_9_LC_5_6_3.C_ON=1'b0;
    defparam beamX_RNII5M_9_LC_5_6_3.SEQ_MODE=4'b0000;
    defparam beamX_RNII5M_9_LC_5_6_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNII5M_9_LC_5_6_3 (
            .in0(N__3124),
            .in1(N__3155),
            .in2(N__3099),
            .in3(N__2834),
            .lcout(),
            .ltout(un18_beamylto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIVEM1_4_LC_5_6_4.C_ON=1'b0;
    defparam beamX_RNIVEM1_4_LC_5_6_4.SEQ_MODE=4'b0000;
    defparam beamX_RNIVEM1_4_LC_5_6_4.LUT_INIT=16'b1101000011000000;
    LogicCell40 beamX_RNIVEM1_4_LC_5_6_4 (
            .in0(N__2660),
            .in1(N__2873),
            .in2(N__2664),
            .in3(N__2906),
            .lcout(un18_beamylt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI8P51_4_LC_5_6_5.C_ON=1'b0;
    defparam beamX_RNI8P51_4_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam beamX_RNI8P51_4_LC_5_6_5.LUT_INIT=16'b0000110100001111;
    LogicCell40 beamX_RNI8P51_4_LC_5_6_5 (
            .in0(N__2907),
            .in1(N__2661),
            .in2(N__2841),
            .in3(N__2874),
            .lcout(un13_beamylt7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNICPU5_10_LC_5_6_7.C_ON=1'b0;
    defparam beamX_RNICPU5_10_LC_5_6_7.SEQ_MODE=4'b0000;
    defparam beamX_RNICPU5_10_LC_5_6_7.LUT_INIT=16'b0001000000000000;
    LogicCell40 beamX_RNICPU5_10_LC_5_6_7 (
            .in0(N__4299),
            .in1(N__2976),
            .in2(N__2915),
            .in3(N__3028),
            .lcout(un3_beamx_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_5_7_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_5_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_5_7_0 (
            .in0(_gnd_net_),
            .in1(N__4352),
            .in2(N__4307),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_RNITP5A_LC_5_7_1.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_RNITP5A_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_RNITP5A_LC_5_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un8_beamx_cry_1_c_RNITP5A_LC_5_7_1 (
            .in0(_gnd_net_),
            .in1(N__2974),
            .in2(_gnd_net_),
            .in3(N__2688),
            .lcout(un8_beamx_cry_1_c_RNITP5AZ0),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_5_7_2.C_ON=1'b1;
    defparam beamX_3_LC_5_7_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_5_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_5_7_2 (
            .in0(_gnd_net_),
            .in1(N__2948),
            .in2(_gnd_net_),
            .in3(N__2685),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__5590),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_5_7_3.C_ON=1'b1;
    defparam beamX_4_LC_5_7_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_5_7_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_5_7_3 (
            .in0(N__4476),
            .in1(N__2911),
            .in2(_gnd_net_),
            .in3(N__2682),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__5590),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_5_7_4.C_ON=1'b1;
    defparam beamX_5_LC_5_7_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_5_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_5_7_4 (
            .in0(_gnd_net_),
            .in1(N__2877),
            .in2(_gnd_net_),
            .in3(N__2679),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__5590),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_5_7_5.C_ON=1'b1;
    defparam beamX_6_LC_5_7_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_5_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_5_7_5 (
            .in0(_gnd_net_),
            .in1(N__2840),
            .in2(_gnd_net_),
            .in3(N__2676),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__5590),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_5_7_6.C_ON=1'b1;
    defparam beamX_7_LC_5_7_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_5_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_5_7_6 (
            .in0(_gnd_net_),
            .in1(N__3159),
            .in2(_gnd_net_),
            .in3(N__2673),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__5590),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_5_7_7.C_ON=1'b1;
    defparam beamX_8_LC_5_7_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_5_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_5_7_7 (
            .in0(_gnd_net_),
            .in1(N__3126),
            .in2(_gnd_net_),
            .in3(N__2670),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__5590),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_5_8_0.C_ON=1'b1;
    defparam beamX_9_LC_5_8_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_5_8_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_5_8_0 (
            .in0(_gnd_net_),
            .in1(N__3094),
            .in2(_gnd_net_),
            .in3(N__2667),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__5589),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_5_8_1.C_ON=1'b0;
    defparam beamX_10_LC_5_8_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_5_8_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_10_LC_5_8_1 (
            .in0(N__4471),
            .in1(N__3022),
            .in2(_gnd_net_),
            .in3(N__2709),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5589),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_5_8_7.C_ON=1'b0;
    defparam beamX_2_LC_5_8_7.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_5_8_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamX_2_LC_5_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3704),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5589),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_1_c_LC_6_2_0.C_ON=1'b1;
    defparam un20_beamy_cry_1_c_LC_6_2_0.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_1_c_LC_6_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un20_beamy_cry_1_c_LC_6_2_0 (
            .in0(_gnd_net_),
            .in1(N__5726),
            .in2(N__3689),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_2_0_),
            .carryout(un20_beamy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_1_c_RNI97C4_LC_6_2_1.C_ON=1'b1;
    defparam un20_beamy_cry_1_c_RNI97C4_LC_6_2_1.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_1_c_RNI97C4_LC_6_2_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un20_beamy_cry_1_c_RNI97C4_LC_6_2_1 (
            .in0(_gnd_net_),
            .in1(N__5345),
            .in2(_gnd_net_),
            .in3(N__2706),
            .lcout(un20_beamy_cry_1_c_RNI97CZ0Z4),
            .ltout(),
            .carryin(un20_beamy_cry_1),
            .carryout(un20_beamy_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_2_c_RNIBAD4_LC_6_2_2.C_ON=1'b1;
    defparam un20_beamy_cry_2_c_RNIBAD4_LC_6_2_2.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_2_c_RNIBAD4_LC_6_2_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un20_beamy_cry_2_c_RNIBAD4_LC_6_2_2 (
            .in0(_gnd_net_),
            .in1(N__4016),
            .in2(_gnd_net_),
            .in3(N__2703),
            .lcout(un20_beamy_cry_2_c_RNIBADZ0Z4),
            .ltout(),
            .carryin(un20_beamy_cry_2),
            .carryout(un20_beamy_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_3_c_RNIDDE4_LC_6_2_3.C_ON=1'b1;
    defparam un20_beamy_cry_3_c_RNIDDE4_LC_6_2_3.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_3_c_RNIDDE4_LC_6_2_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 un20_beamy_cry_3_c_RNIDDE4_LC_6_2_3 (
            .in0(_gnd_net_),
            .in1(N__4176),
            .in2(_gnd_net_),
            .in3(N__2700),
            .lcout(un20_beamy_cry_3_c_RNIDDEZ0Z4),
            .ltout(),
            .carryin(un20_beamy_cry_3),
            .carryout(un20_beamy_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_4_c_RNIFGF4_LC_6_2_4.C_ON=1'b1;
    defparam un20_beamy_cry_4_c_RNIFGF4_LC_6_2_4.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_4_c_RNIFGF4_LC_6_2_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un20_beamy_cry_4_c_RNIFGF4_LC_6_2_4 (
            .in0(_gnd_net_),
            .in1(N__3957),
            .in2(_gnd_net_),
            .in3(N__2697),
            .lcout(un20_beamy_cry_4_c_RNIFGFZ0Z4),
            .ltout(),
            .carryin(un20_beamy_cry_4),
            .carryout(un20_beamy_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_5_c_RNIHJG4_LC_6_2_5.C_ON=1'b1;
    defparam un20_beamy_cry_5_c_RNIHJG4_LC_6_2_5.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_5_c_RNIHJG4_LC_6_2_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un20_beamy_cry_5_c_RNIHJG4_LC_6_2_5 (
            .in0(_gnd_net_),
            .in1(N__4556),
            .in2(_gnd_net_),
            .in3(N__2694),
            .lcout(un20_beamy_cry_5_c_RNIHJGZ0Z4),
            .ltout(),
            .carryin(un20_beamy_cry_5),
            .carryout(un20_beamy_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un20_beamy_cry_6_c_RNIJMH4_LC_6_2_6.C_ON=1'b1;
    defparam un20_beamy_cry_6_c_RNIJMH4_LC_6_2_6.SEQ_MODE=4'b0000;
    defparam un20_beamy_cry_6_c_RNIJMH4_LC_6_2_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 un20_beamy_cry_6_c_RNIJMH4_LC_6_2_6 (
            .in0(_gnd_net_),
            .in1(N__4068),
            .in2(_gnd_net_),
            .in3(N__2691),
            .lcout(un20_beamy_cry_6_c_RNIJMHZ0Z4),
            .ltout(),
            .carryin(un20_beamy_cry_6),
            .carryout(un20_beamy_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_8_LC_6_2_7.C_ON=1'b1;
    defparam beamY_8_LC_6_2_7.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_6_2_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_6_2_7 (
            .in0(_gnd_net_),
            .in1(N__4123),
            .in2(_gnd_net_),
            .in3(N__2739),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un20_beamy_cry_7),
            .carryout(un20_beamy_cry_8),
            .clk(N__5597),
            .ce(N__4467),
            .sr(_gnd_net_));
    defparam beamY_9_LC_6_3_0.C_ON=1'b0;
    defparam beamY_9_LC_6_3_0.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_6_3_0.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamY_9_LC_6_3_0 (
            .in0(N__3902),
            .in1(N__3191),
            .in2(_gnd_net_),
            .in3(N__2736),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5595),
            .ce(N__4468),
            .sr(_gnd_net_));
    defparam beamY_RNID825_6_LC_6_4_0.C_ON=1'b0;
    defparam beamY_RNID825_6_LC_6_4_0.SEQ_MODE=4'b0000;
    defparam beamY_RNID825_6_LC_6_4_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 beamY_RNID825_6_LC_6_4_0 (
            .in0(N__2721),
            .in1(N__4560),
            .in2(_gnd_net_),
            .in3(N__4134),
            .lcout(),
            .ltout(un5_beamx_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DLC_5_LC_6_4_1.C_ON=1'b0;
    defparam beamY_RNI9DLC_5_LC_6_4_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DLC_5_LC_6_4_1.LUT_INIT=16'b0000000001000000;
    LogicCell40 beamY_RNI9DLC_5_LC_6_4_1 (
            .in0(N__5352),
            .in1(N__2727),
            .in2(N__2733),
            .in3(N__3953),
            .lcout(beamY_RNI9DLCZ0Z_5),
            .ltout(beamY_RNI9DLCZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_6_4_2.C_ON=1'b0;
    defparam beamY_0_LC_6_4_2.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_6_4_2.LUT_INIT=16'b0000001111001100;
    LogicCell40 beamY_0_LC_6_4_2 (
            .in0(_gnd_net_),
            .in1(N__3677),
            .in2(N__2730),
            .in3(N__4457),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5594),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9425_0_LC_6_4_3.C_ON=1'b0;
    defparam beamY_RNI9425_0_LC_6_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI9425_0_LC_6_4_3.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_RNI9425_0_LC_6_4_3 (
            .in0(N__5713),
            .in1(N__3888),
            .in2(N__3685),
            .in3(N__4066),
            .lcout(un5_beamx_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIJ0H2_4_LC_6_4_4.C_ON=1'b0;
    defparam beamY_RNIJ0H2_4_LC_6_4_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIJ0H2_4_LC_6_4_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 beamY_RNIJ0H2_4_LC_6_4_4 (
            .in0(_gnd_net_),
            .in1(N__4169),
            .in2(_gnd_net_),
            .in3(N__4015),
            .lcout(un5_beamx_2),
            .ltout(un5_beamx_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI5NA6_5_LC_6_4_5.C_ON=1'b0;
    defparam beamY_RNI5NA6_5_LC_6_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI5NA6_5_LC_6_4_5.LUT_INIT=16'b0000000000010011;
    LogicCell40 beamY_RNI5NA6_5_LC_6_4_5 (
            .in0(N__5351),
            .in1(N__3887),
            .in2(N__2715),
            .in3(N__3952),
            .lcout(),
            .ltout(un8_beamylto9_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_6_LC_6_4_6.C_ON=1'b0;
    defparam beamY_RNISI4A_6_LC_6_4_6.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_6_LC_6_4_6.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamY_RNISI4A_6_LC_6_4_6 (
            .in0(N__4065),
            .in1(N__4559),
            .in2(N__2712),
            .in3(N__4133),
            .lcout(un8_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_0_3_LC_6_5_0.C_ON=1'b0;
    defparam beamY_RNIHUG2_0_3_LC_6_5_0.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_0_3_LC_6_5_0.LUT_INIT=16'b0000000001010101;
    LogicCell40 beamY_RNIHUG2_0_3_LC_6_5_0 (
            .in0(N__4020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5346),
            .lcout(),
            .ltout(un4_beamylt6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_4_LC_6_5_1.C_ON=1'b0;
    defparam beamY_RNI2KA6_4_LC_6_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_4_LC_6_5_1.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_RNI2KA6_4_LC_6_5_1 (
            .in0(N__4180),
            .in1(N__3961),
            .in2(N__2802),
            .in3(N__4557),
            .lcout(),
            .ltout(un4_beamylt8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_7_LC_6_5_2.C_ON=1'b0;
    defparam beamY_RNISI4A_7_LC_6_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_7_LC_6_5_2.LUT_INIT=16'b1100110011001000;
    LogicCell40 beamY_RNISI4A_7_LC_6_5_2 (
            .in0(N__4077),
            .in1(N__3903),
            .in2(N__2799),
            .in3(N__4135),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_6_5_4.C_ON=1'b0;
    defparam beamY_1_LC_6_5_4.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_6_5_4.LUT_INIT=16'b0101001001110000;
    LogicCell40 beamY_1_LC_6_5_4 (
            .in0(N__4446),
            .in1(N__3192),
            .in2(N__5730),
            .in3(N__3681),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5593),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIKVE6_3_LC_6_6_0.C_ON=1'b0;
    defparam beamX_RNIKVE6_3_LC_6_6_0.SEQ_MODE=4'b0000;
    defparam beamX_RNIKVE6_3_LC_6_6_0.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamX_RNIKVE6_3_LC_6_6_0 (
            .in0(N__2838),
            .in1(N__2946),
            .in2(N__2796),
            .in3(N__4358),
            .lcout(),
            .ltout(un3_beamx_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI5457_5_LC_6_6_1.C_ON=1'b0;
    defparam beamX_RNI5457_5_LC_6_6_1.SEQ_MODE=4'b0000;
    defparam beamX_RNI5457_5_LC_6_6_1.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNI5457_5_LC_6_6_1 (
            .in0(N__2999),
            .in1(N__3157),
            .in2(N__2787),
            .in3(N__2875),
            .lcout(beamX_RNI5457Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_RNO_0_LC_6_6_3.C_ON=1'b0;
    defparam HSync_1_RNO_0_LC_6_6_3.SEQ_MODE=4'b0000;
    defparam HSync_1_RNO_0_LC_6_6_3.LUT_INIT=16'b1000000000000000;
    LogicCell40 HSync_1_RNO_0_LC_6_6_3 (
            .in0(N__2947),
            .in1(N__2876),
            .in2(N__2916),
            .in3(N__2839),
            .lcout(),
            .ltout(un1_beamxlt10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_6_6_4.C_ON=1'b0;
    defparam HSync_1_LC_6_6_4.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_6_6_4.LUT_INIT=16'b1111111011111111;
    LogicCell40 HSync_1_LC_6_6_4 (
            .in0(N__3158),
            .in1(N__3030),
            .in2(N__2784),
            .in3(N__3000),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5592),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIR4B_9_LC_6_6_5.C_ON=1'b0;
    defparam beamX_RNIR4B_9_LC_6_6_5.SEQ_MODE=4'b0000;
    defparam beamX_RNIR4B_9_LC_6_6_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_RNIR4B_9_LC_6_6_5 (
            .in0(_gnd_net_),
            .in1(N__3098),
            .in2(_gnd_net_),
            .in3(N__3125),
            .lcout(un1_beamx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIT9ER_10_LC_6_6_6.C_ON=1'b0;
    defparam beamX_RNIT9ER_10_LC_6_6_6.SEQ_MODE=4'b0000;
    defparam beamX_RNIT9ER_10_LC_6_6_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamX_RNIT9ER_10_LC_6_6_6 (
            .in0(N__2745),
            .in1(N__3048),
            .in2(N__3039),
            .in3(N__3029),
            .lcout(),
            .ltout(un15_beamy_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNISO4T_7_LC_6_6_7.C_ON=1'b0;
    defparam beamX_RNISO4T_7_LC_6_6_7.SEQ_MODE=4'b0000;
    defparam beamX_RNISO4T_7_LC_6_6_7.LUT_INIT=16'b0111000001010000;
    LogicCell40 beamX_RNISO4T_7_LC_6_6_7 (
            .in0(N__2998),
            .in1(N__2988),
            .in2(N__2982),
            .in3(N__3156),
            .lcout(un15_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_0_c_LC_6_7_0.C_ON=1'b1;
    defparam un5_visiblex_1_cry_0_c_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_0_c_LC_6_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_visiblex_1_cry_0_c_LC_6_7_0 (
            .in0(_gnd_net_),
            .in1(N__4337),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(un5_visiblex_1_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_0_c_RNI1IJC_LC_6_7_1.C_ON=1'b1;
    defparam un5_visiblex_1_cry_0_c_RNI1IJC_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_0_c_RNI1IJC_LC_6_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_1_cry_0_c_RNI1IJC_LC_6_7_1 (
            .in0(_gnd_net_),
            .in1(N__4297),
            .in2(_gnd_net_),
            .in3(N__2979),
            .lcout(un5_visiblex_1_n_31),
            .ltout(),
            .carryin(un5_visiblex_1_cry_0),
            .carryout(un5_visiblex_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_1_c_RNI3LKC_LC_6_7_2.C_ON=1'b1;
    defparam un5_visiblex_1_cry_1_c_RNI3LKC_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_1_c_RNI3LKC_LC_6_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_1_cry_1_c_RNI3LKC_LC_6_7_2 (
            .in0(_gnd_net_),
            .in1(N__2968),
            .in2(_gnd_net_),
            .in3(N__2952),
            .lcout(un5_visiblex_1_n_30),
            .ltout(),
            .carryin(un5_visiblex_1_cry_1),
            .carryout(un5_visiblex_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_2_c_RNI5OLC_LC_6_7_3.C_ON=1'b1;
    defparam un5_visiblex_1_cry_2_c_RNI5OLC_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_2_c_RNI5OLC_LC_6_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_1_cry_2_c_RNI5OLC_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(N__2942),
            .in2(N__5458),
            .in3(N__2919),
            .lcout(un1_visiblex_24),
            .ltout(),
            .carryin(un5_visiblex_1_cry_2),
            .carryout(un5_visiblex_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_3_c_RNI7RMC_LC_6_7_4.C_ON=1'b1;
    defparam un5_visiblex_1_cry_3_c_RNI7RMC_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_3_c_RNI7RMC_LC_6_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_1_cry_3_c_RNI7RMC_LC_6_7_4 (
            .in0(_gnd_net_),
            .in1(N__2905),
            .in2(_gnd_net_),
            .in3(N__2880),
            .lcout(un5_visiblex_1_n_28),
            .ltout(),
            .carryin(un5_visiblex_1_cry_3),
            .carryout(un5_visiblex_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_4_c_RNI9UNC_LC_6_7_5.C_ON=1'b1;
    defparam un5_visiblex_1_cry_4_c_RNI9UNC_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_4_c_RNI9UNC_LC_6_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_1_cry_4_c_RNI9UNC_LC_6_7_5 (
            .in0(_gnd_net_),
            .in1(N__2872),
            .in2(_gnd_net_),
            .in3(N__2844),
            .lcout(un5_visiblex_1_n_27),
            .ltout(),
            .carryin(un5_visiblex_1_cry_4),
            .carryout(un5_visiblex_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_5_c_RNIB1PC_LC_6_7_6.C_ON=1'b1;
    defparam un5_visiblex_1_cry_5_c_RNIB1PC_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_5_c_RNIB1PC_LC_6_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_1_cry_5_c_RNIB1PC_LC_6_7_6 (
            .in0(_gnd_net_),
            .in1(N__2833),
            .in2(N__5459),
            .in3(N__2805),
            .lcout(un5_visiblex_1_n_26),
            .ltout(),
            .carryin(un5_visiblex_1_cry_5),
            .carryout(un5_visiblex_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_6_c_RNID4QC_LC_6_7_7.C_ON=1'b1;
    defparam un5_visiblex_1_cry_6_c_RNID4QC_LC_6_7_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_6_c_RNID4QC_LC_6_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_visiblex_1_cry_6_c_RNID4QC_LC_6_7_7 (
            .in0(_gnd_net_),
            .in1(N__3154),
            .in2(_gnd_net_),
            .in3(N__3129),
            .lcout(un5_visiblex_1_n_25),
            .ltout(),
            .carryin(un5_visiblex_1_cry_6),
            .carryout(un5_visiblex_1_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_7_c_RNIF7RC_LC_6_8_0.C_ON=1'b1;
    defparam un5_visiblex_1_cry_7_c_RNIF7RC_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_7_c_RNIF7RC_LC_6_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_visiblex_1_cry_7_c_RNIF7RC_LC_6_8_0 (
            .in0(_gnd_net_),
            .in1(N__3123),
            .in2(N__5460),
            .in3(N__3102),
            .lcout(un5_visiblex_1_n_24),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(un5_visiblex_1_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_8_c_RNIHASC_LC_6_8_1.C_ON=1'b0;
    defparam un5_visiblex_1_cry_8_c_RNIHASC_LC_6_8_1.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_8_c_RNIHASC_LC_6_8_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_visiblex_1_cry_8_c_RNIHASC_LC_6_8_1 (
            .in0(_gnd_net_),
            .in1(N__3087),
            .in2(_gnd_net_),
            .in3(N__3066),
            .lcout(un5_visiblex_1_n_23),
            .ltout(un5_visiblex_1_n_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_8_c_RNIHASC_1_LC_6_8_2.C_ON=1'b0;
    defparam un5_visiblex_1_cry_8_c_RNIHASC_1_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_8_c_RNIHASC_1_LC_6_8_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 un5_visiblex_1_cry_8_c_RNIHASC_1_LC_6_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3063),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_s_5_sf),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_LC_7_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3594),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_7_2_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_7_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_7_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3I151_LC_7_2_1 (
            .in0(_gnd_net_),
            .in1(N__5411),
            .in2(N__3231),
            .in3(N__3060),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNI3IZ0Z151),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_7_2_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_7_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_7_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4K251_LC_7_2_2 (
            .in0(_gnd_net_),
            .in1(N__3720),
            .in2(N__5442),
            .in3(N__3057),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3_c_RNI4KZ0Z251),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_7_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3054),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_7_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3051),
            .in3(N__4663),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIGR79_7_LC_7_2_6.C_ON=1'b0;
    defparam beamY_fast_RNIGR79_7_LC_7_2_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIGR79_7_LC_7_2_6.LUT_INIT=16'b1111111111111010;
    LogicCell40 beamY_fast_RNIGR79_7_LC_7_2_6 (
            .in0(N__4102),
            .in1(_gnd_net_),
            .in2(N__3585),
            .in3(N__3567),
            .lcout(beamY_fast_RNIGR79Z0Z_7),
            .ltout(beamY_fast_RNIGR79Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIALEQ_0_9_LC_7_2_7.C_ON=1'b0;
    defparam beamY_RNIALEQ_0_9_LC_7_2_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIALEQ_0_9_LC_7_2_7.LUT_INIT=16'b0011110000110011;
    LogicCell40 beamY_RNIALEQ_0_9_LC_7_2_7 (
            .in0(_gnd_net_),
            .in1(N__3886),
            .in2(N__3234),
            .in3(N__3644),
            .lcout(beamY_RNIALEQ_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_3_LC_7_3_0.C_ON=1'b0;
    defparam beamY_3_LC_7_3_0.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_7_3_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_3_LC_7_3_0 (
            .in0(_gnd_net_),
            .in1(N__3221),
            .in2(_gnd_net_),
            .in3(N__3185),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam beamY_fast_7_LC_7_3_1.C_ON=1'b0;
    defparam beamY_fast_7_LC_7_3_1.SEQ_MODE=4'b1000;
    defparam beamY_fast_7_LC_7_3_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_fast_7_LC_7_3_1 (
            .in0(N__3190),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3204),
            .lcout(beamY_fastZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam beamY_fast_4_LC_7_3_2.C_ON=1'b0;
    defparam beamY_fast_4_LC_7_3_2.SEQ_MODE=4'b1000;
    defparam beamY_fast_4_LC_7_3_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 beamY_fast_4_LC_7_3_2 (
            .in0(N__3213),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3189),
            .lcout(beamY_fastZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam beamY_5_LC_7_3_3.C_ON=1'b0;
    defparam beamY_5_LC_7_3_3.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_7_3_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_5_LC_7_3_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3272),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam beamY_fast_3_LC_7_3_4.C_ON=1'b0;
    defparam beamY_fast_3_LC_7_3_4.SEQ_MODE=4'b1000;
    defparam beamY_fast_3_LC_7_3_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_fast_3_LC_7_3_4 (
            .in0(_gnd_net_),
            .in1(N__3222),
            .in2(_gnd_net_),
            .in3(N__3188),
            .lcout(beamY_fastZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam beamY_4_LC_7_3_5.C_ON=1'b0;
    defparam beamY_4_LC_7_3_5.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_7_3_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 beamY_4_LC_7_3_5 (
            .in0(N__3186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3212),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam beamY_7_LC_7_3_6.C_ON=1'b0;
    defparam beamY_7_LC_7_3_6.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_7_3_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 beamY_7_LC_7_3_6 (
            .in0(_gnd_net_),
            .in1(N__3203),
            .in2(_gnd_net_),
            .in3(N__3187),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam beamY_fast_5_LC_7_3_7.C_ON=1'b0;
    defparam beamY_fast_5_LC_7_3_7.SEQ_MODE=4'b1000;
    defparam beamY_fast_5_LC_7_3_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_5_LC_7_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3273),
            .lcout(beamY_fastZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5598),
            .ce(N__4469),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_4_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_4_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_4_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_16_LC_7_5_0.C_ON=1'b0;
    defparam Pixel_1_RNO_16_LC_7_5_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_16_LC_7_5_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 Pixel_1_RNO_16_LC_7_5_0 (
            .in0(_gnd_net_),
            .in1(N__4022),
            .in2(_gnd_net_),
            .in3(N__5348),
            .lcout(un12_visiblexlt9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_4_LC_7_5_2.C_ON=1'b0;
    defparam Pixel_1_RNO_4_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_4_LC_7_5_2.LUT_INIT=16'b0010100000000000;
    LogicCell40 Pixel_1_RNO_4_LC_7_5_2 (
            .in0(N__3264),
            .in1(N__3904),
            .in2(N__3633),
            .in3(N__3336),
            .lcout(un13_visiblex_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI8CP3_1_LC_7_5_4.C_ON=1'b0;
    defparam beamY_RNI8CP3_1_LC_7_5_4.SEQ_MODE=4'b0000;
    defparam beamY_RNI8CP3_1_LC_7_5_4.LUT_INIT=16'b0010001011001100;
    LogicCell40 beamY_RNI8CP3_1_LC_7_5_4 (
            .in0(N__5703),
            .in1(N__4021),
            .in2(_gnd_net_),
            .in3(N__5347),
            .lcout(font_un7_pixellt9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_RNO_0_LC_7_5_6.C_ON=1'b0;
    defparam VSync_1_RNO_0_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam VSync_1_RNO_0_LC_7_5_6.LUT_INIT=16'b0001000100110011;
    LogicCell40 VSync_1_RNO_0_LC_7_5_6 (
            .in0(N__5704),
            .in1(N__4181),
            .in2(_gnd_net_),
            .in3(N__5349),
            .lcout(un1_beamylto9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_11_LC_7_6_0.C_ON=1'b0;
    defparam Pixel_1_RNO_11_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_11_LC_7_6_0.LUT_INIT=16'b0000000000010000;
    LogicCell40 Pixel_1_RNO_11_LC_7_6_0 (
            .in0(N__4262),
            .in1(N__3814),
            .in2(N__3252),
            .in3(N__3509),
            .lcout(un13_visiblex_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_15_LC_7_6_1.C_ON=1'b0;
    defparam Pixel_1_RNO_15_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_15_LC_7_6_1.LUT_INIT=16'b0001000100010011;
    LogicCell40 Pixel_1_RNO_15_LC_7_6_1 (
            .in0(N__5140),
            .in1(N__3258),
            .in2(N__3321),
            .in3(N__3306),
            .lcout(un13_visiblex_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIU8361_0_LC_7_6_2.C_ON=1'b0;
    defparam beamX_RNIU8361_0_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam beamX_RNIU8361_0_LC_7_6_2.LUT_INIT=16'b1100110010001100;
    LogicCell40 beamX_RNIU8361_0_LC_7_6_2 (
            .in0(N__3304),
            .in1(N__5136),
            .in2(N__4359),
            .in3(N__3316),
            .lcout(),
            .ltout(font_un14_pixellt9_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIUQF32_0_LC_7_6_3.C_ON=1'b0;
    defparam beamX_RNIUQF32_0_LC_7_6_3.SEQ_MODE=4'b0000;
    defparam beamX_RNIUQF32_0_LC_7_6_3.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamX_RNIUQF32_0_LC_7_6_3 (
            .in0(N__3243),
            .in1(N__3813),
            .in2(N__3237),
            .in3(N__4261),
            .lcout(Pixel_0_sqmuxa_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_4_c_RNIAG3A1_LC_7_6_5.C_ON=1'b0;
    defparam un5_visiblex_1_cry_4_c_RNIAG3A1_LC_7_6_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_4_c_RNIAG3A1_LC_7_6_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 un5_visiblex_1_cry_4_c_RNIAG3A1_LC_7_6_5 (
            .in0(N__5485),
            .in1(N__5231),
            .in2(N__5092),
            .in3(N__3432),
            .lcout(un13_visiblex_5),
            .ltout(un13_visiblex_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNINUI05_0_LC_7_6_6.C_ON=1'b0;
    defparam beamX_RNINUI05_0_LC_7_6_6.SEQ_MODE=4'b0000;
    defparam beamX_RNINUI05_0_LC_7_6_6.LUT_INIT=16'b0000000001000000;
    LogicCell40 beamX_RNINUI05_0_LC_7_6_6 (
            .in0(N__3294),
            .in1(N__3330),
            .in2(N__3324),
            .in3(N__3510),
            .lcout(Pixel_0_sqmuxa_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIU8361_0_0_LC_7_6_7.C_ON=1'b0;
    defparam beamX_RNIU8361_0_0_LC_7_6_7.SEQ_MODE=4'b0000;
    defparam beamX_RNIU8361_0_0_LC_7_6_7.LUT_INIT=16'b0000000000000100;
    LogicCell40 beamX_RNIU8361_0_0_LC_7_6_7 (
            .in0(N__3317),
            .in1(N__4356),
            .in2(N__5144),
            .in3(N__3305),
            .lcout(N_159),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_7_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_LC_7_7_0 (
            .in0(_gnd_net_),
            .in1(N__4257),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKV_LC_7_7_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKV_LC_7_7_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKV_LC_7_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKV_LC_7_7_1 (
            .in0(_gnd_net_),
            .in1(N__3366),
            .in2(N__3441),
            .in3(N__3288),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4_c_RNI0SKVZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUD1_LC_7_7_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUD1_LC_7_7_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUD1_LC_7_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUD1_LC_7_7_2 (
            .in0(_gnd_net_),
            .in1(N__3356),
            .in2(N__3405),
            .in3(N__3285),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5_c_RNIRJUDZ0Z1),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISJ3S2_LC_7_7_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISJ3S2_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISJ3S2_LC_7_7_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6_c_RNISJ3S2_LC_7_7_3 (
            .in0(N__3788),
            .in1(N__3342),
            .in2(N__3393),
            .in3(N__3282),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_LC_7_7_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_LC_7_7_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_LC_7_7_4 (
            .in0(N__3357),
            .in1(N__3503),
            .in2(N__3381),
            .in3(N__3279),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1),
            .ltout(un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2EZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_0_LC_7_7_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_0_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_0_LC_7_7_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un54_sum_cry_7_c_RNIVR2E1_0_LC_7_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3276),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_7_c_RNIF7RC_0_LC_7_7_6.C_ON=1'b0;
    defparam un5_visiblex_1_cry_7_c_RNIF7RC_0_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_7_c_RNIF7RC_0_LC_7_7_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_1_cry_7_c_RNIF7RC_0_LC_7_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3428),
            .lcout(un5_visiblex_1_n_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_8_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__3427),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3R_LC_7_8_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3R_LC_7_8_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3R_LC_7_8_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3R_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__3411),
            .in2(_gnd_net_),
            .in3(N__3396),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4_c_RNI9T3RZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4R_LC_7_8_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4R_LC_7_8_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4R_LC_7_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4R_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(N__3483),
            .in2(N__5443),
            .in3(N__3384),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5_c_RNIAV4RZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_7_8_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_7_8_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_7_8_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_LUT4_0_LC_7_8_3 (
            .in0(_gnd_net_),
            .in1(N__3502),
            .in2(_gnd_net_),
            .in3(N__3372),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_7_8_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_7_8_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_7_8_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_LUT4_0_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3369),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO),
            .ltout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_7_8_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_7_8_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_7_8_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_LC_7_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3360),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0),
            .ltout(un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAEZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_7_8_6.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_7_8_6.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_7_8_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un47_sum_cry_7_c_RNIROAE_0_LC_7_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3345),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_8_c_RNIHASC_0_LC_7_8_7.C_ON=1'b0;
    defparam un5_visiblex_1_cry_8_c_RNIHASC_0_LC_7_8_7.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_8_c_RNIHASC_0_LC_7_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_1_cry_8_c_RNIHASC_0_LC_7_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3501),
            .lcout(un5_visiblex_1_cry_8_c_RNIHASCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_1_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_LC_8_1_0 (
            .in0(_gnd_net_),
            .in1(N__4609),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250Q_LC_8_1_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250Q_LC_8_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250Q_LC_8_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250Q_LC_8_1_1 (
            .in0(_gnd_net_),
            .in1(N__3525),
            .in2(N__5447),
            .in3(N__3477),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2_c_RNI250QZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_1_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPS51_LC_8_1_2 (
            .in0(_gnd_net_),
            .in1(N__3474),
            .in2(N__5449),
            .in3(N__3468),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3_c_RNIRPSZ0Z51),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_1_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTU51_LC_8_1_3 (
            .in0(_gnd_net_),
            .in1(N__3465),
            .in2(N__5448),
            .in3(N__3459),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNITTUZ0Z51),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_1_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_1_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_8_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4664),
            .in3(N__3456),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_1_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJB_LC_8_1_5 (
            .in0(_gnd_net_),
            .in1(N__3453),
            .in2(_gnd_net_),
            .in3(N__3447),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_6_c_RNIMEJBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIH1_LC_8_1_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIH1_LC_8_1_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIH1_LC_8_1_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIH1_LC_8_1_6 (
            .in0(N__4698),
            .in1(_gnd_net_),
            .in2(N__3444),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_cry_4_c_RNIJCIHZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIIGUB_2_LC_8_2_0.C_ON=1'b0;
    defparam beamY_fast_RNIIGUB_2_LC_8_2_0.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIIGUB_2_LC_8_2_0.LUT_INIT=16'b1010000000000000;
    LogicCell40 beamY_fast_RNIIGUB_2_LC_8_2_0 (
            .in0(N__4491),
            .in1(_gnd_net_),
            .in2(N__3750),
            .in3(N__3765),
            .lcout(un5_visibley_c3),
            .ltout(un5_visibley_c3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIJ9FI_5_LC_8_2_1.C_ON=1'b0;
    defparam beamY_fast_RNIJ9FI_5_LC_8_2_1.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIJ9FI_5_LC_8_2_1.LUT_INIT=16'b1100110011001001;
    LogicCell40 beamY_fast_RNIJ9FI_5_LC_8_2_1 (
            .in0(N__3566),
            .in1(N__4076),
            .in2(N__3600),
            .in3(N__4532),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_0_LC_8_2_2.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_0_LC_8_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_0_LC_8_2_2.LUT_INIT=16'b1111000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_0_LC_8_2_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3749),
            .in3(N__3764),
            .lcout(),
            .ltout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_8_2_3.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_8_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_8_2_3.LUT_INIT=16'b1010101010010101;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNO_LC_8_2_3 (
            .in0(N__4124),
            .in1(N__4490),
            .in2(N__3597),
            .in3(N__3551),
            .lcout(un1_beamY_if_generate_plus_mult1_un33_sum_cry_2_c_RNOZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIU8LB1_8_LC_8_2_4.C_ON=1'b0;
    defparam beamY_RNIU8LB1_8_LC_8_2_4.SEQ_MODE=4'b0000;
    defparam beamY_RNIU8LB1_8_LC_8_2_4.LUT_INIT=16'b0000000100110010;
    LogicCell40 beamY_RNIU8LB1_8_LC_8_2_4 (
            .in0(N__3552),
            .in1(N__4611),
            .in2(N__3540),
            .in3(N__4126),
            .lcout(un13_visiblex_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9LFE_6_LC_8_2_5.C_ON=1'b0;
    defparam beamY_RNI9LFE_6_LC_8_2_5.SEQ_MODE=4'b0000;
    defparam beamY_RNI9LFE_6_LC_8_2_5.LUT_INIT=16'b1100110010011001;
    LogicCell40 beamY_RNI9LFE_6_LC_8_2_5 (
            .in0(N__3947),
            .in1(N__4533),
            .in2(_gnd_net_),
            .in3(N__3536),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIRPUB_6_LC_8_2_6.C_ON=1'b0;
    defparam beamY_fast_RNIRPUB_6_LC_8_2_6.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIRPUB_6_LC_8_2_6.LUT_INIT=16'b1111111111111100;
    LogicCell40 beamY_fast_RNIRPUB_6_LC_8_2_6 (
            .in0(_gnd_net_),
            .in1(N__4583),
            .in2(N__3584),
            .in3(N__3565),
            .lcout(un5_visibley_c6_0_0_0),
            .ltout(un5_visibley_c6_0_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBV5P_8_LC_8_2_7.C_ON=1'b0;
    defparam beamY_RNIBV5P_8_LC_8_2_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIBV5P_8_LC_8_2_7.LUT_INIT=16'b0101010101011010;
    LogicCell40 beamY_RNIBV5P_8_LC_8_2_7 (
            .in0(N__4125),
            .in1(_gnd_net_),
            .in2(N__3543),
            .in3(N__3535),
            .lcout(beamY_RNIBV5PZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI6125_4_LC_8_3_0.C_ON=1'b0;
    defparam beamY_RNI6125_4_LC_8_3_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI6125_4_LC_8_3_0.LUT_INIT=16'b1000000001111111;
    LogicCell40 beamY_RNI6125_4_LC_8_3_0 (
            .in0(N__4004),
            .in1(N__5306),
            .in2(N__4182),
            .in3(N__3948),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum),
            .ltout(un1_beamY_if_generate_plus_mult1_un54_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIDV6V1_8_LC_8_3_1.C_ON=1'b0;
    defparam beamY_RNIDV6V1_8_LC_8_3_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIDV6V1_8_LC_8_3_1.LUT_INIT=16'b0000000000001010;
    LogicCell40 beamY_RNIDV6V1_8_LC_8_3_1 (
            .in0(N__3519),
            .in1(_gnd_net_),
            .in2(N__3513),
            .in3(N__4846),
            .lcout(Pixel_0_sqmuxa_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_RNIR3UF_6_LC_8_3_2.C_ON=1'b0;
    defparam beamY_fast_RNIR3UF_6_LC_8_3_2.SEQ_MODE=4'b0000;
    defparam beamY_fast_RNIR3UF_6_LC_8_3_2.LUT_INIT=16'b0000011100001111;
    LogicCell40 beamY_fast_RNIR3UF_6_LC_8_3_2 (
            .in0(N__3763),
            .in1(N__3742),
            .in2(N__4587),
            .in3(N__4489),
            .lcout(un5_visibley_ac0_11_0_1),
            .ltout(un5_visibley_ac0_11_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIALEQ_9_LC_8_3_3.C_ON=1'b0;
    defparam beamY_RNIALEQ_9_LC_8_3_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIALEQ_9_LC_8_3_3.LUT_INIT=16'b1100110000111100;
    LogicCell40 beamY_RNIALEQ_9_LC_8_3_3 (
            .in0(_gnd_net_),
            .in1(N__3895),
            .in2(N__3729),
            .in3(N__3726),
            .lcout(beamY_RNIALEQZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_8_3_5.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_8_3_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_8_3_5.LUT_INIT=16'b0110011001100110;
    LogicCell40 beamY_RNIHUG2_3_LC_8_3_5 (
            .in0(N__5307),
            .in1(N__4005),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum),
            .ltout(un1_beamY_if_generate_plus_mult1_un68_sum_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI0R15_1_LC_8_3_6.C_ON=1'b0;
    defparam beamY_RNI0R15_1_LC_8_3_6.SEQ_MODE=4'b0000;
    defparam beamY_RNI0R15_1_LC_8_3_6.LUT_INIT=16'b0000001100000000;
    LogicCell40 beamY_RNI0R15_1_LC_8_3_6 (
            .in0(_gnd_net_),
            .in1(N__5731),
            .in2(N__3714),
            .in3(N__5308),
            .lcout(),
            .ltout(font_un11_pixellto9_7_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIQ0DS_1_LC_8_3_7.C_ON=1'b0;
    defparam beamY_RNIQ0DS_1_LC_8_3_7.SEQ_MODE=4'b0000;
    defparam beamY_RNIQ0DS_1_LC_8_3_7.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamY_RNIQ0DS_1_LC_8_3_7 (
            .in0(N__5220),
            .in1(N__5183),
            .in2(N__3711),
            .in3(N__4845),
            .lcout(font_un11_pixel_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_5_LC_8_4_0.C_ON=1'b0;
    defparam Pixel_1_RNO_5_LC_8_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_5_LC_8_4_0.LUT_INIT=16'b1011000010111011;
    LogicCell40 Pixel_1_RNO_5_LC_8_4_0 (
            .in0(N__3708),
            .in1(N__4272),
            .in2(N__3690),
            .in3(N__5818),
            .lcout(),
            .ltout(font_un26_pixel_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_1_LC_8_4_1.C_ON=1'b0;
    defparam Pixel_1_RNO_1_LC_8_4_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_1_LC_8_4_1.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_1_RNO_1_LC_8_4_1 (
            .in0(N__4206),
            .in1(N__4215),
            .in2(N__3648),
            .in3(N__3606),
            .lcout(d_N_3_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUNJ_7_LC_8_4_2.C_ON=1'b0;
    defparam beamY_RNIHUNJ_7_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUNJ_7_LC_8_4_2.LUT_INIT=16'b1111111111111011;
    LogicCell40 beamY_RNIHUNJ_7_LC_8_4_2 (
            .in0(N__4067),
            .in1(N__3645),
            .in2(N__3962),
            .in3(N__4136),
            .lcout(un5_visibley_c7),
            .ltout(un5_visibley_c7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI1K0I6_9_LC_8_4_3.C_ON=1'b0;
    defparam beamY_RNI1K0I6_9_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNI1K0I6_9_LC_8_4_3.LUT_INIT=16'b0000001000100000;
    LogicCell40 beamY_RNI1K0I6_9_LC_8_4_3 (
            .in0(N__3624),
            .in1(N__3615),
            .in2(N__3609),
            .in3(N__3905),
            .lcout(Pixel_0_sqmuxa_7),
            .ltout(Pixel_0_sqmuxa_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_0_LC_8_4_4.C_ON=1'b0;
    defparam Pixel_1_RNO_0_LC_8_4_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_0_LC_8_4_4.LUT_INIT=16'b0100010001001100;
    LogicCell40 Pixel_1_RNO_0_LC_8_4_4 (
            .in0(N__4214),
            .in1(N__4205),
            .in2(N__4191),
            .in3(N__4188),
            .lcout(Pixel_5_N_3_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIBFP3_4_LC_8_4_5.C_ON=1'b0;
    defparam beamY_RNIBFP3_4_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIBFP3_4_LC_8_4_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 beamY_RNIBFP3_4_LC_8_4_5 (
            .in0(N__5326),
            .in1(N__4168),
            .in2(_gnd_net_),
            .in3(N__4006),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_RNO_1_LC_8_5_4.C_ON=1'b0;
    defparam VSync_1_RNO_1_LC_8_5_4.SEQ_MODE=4'b0000;
    defparam VSync_1_RNO_1_LC_8_5_4.LUT_INIT=16'b0000000000000001;
    LogicCell40 VSync_1_RNO_1_LC_8_5_4 (
            .in0(N__4137),
            .in1(N__4072),
            .in2(N__4026),
            .in3(N__4558),
            .lcout(),
            .ltout(un1_beamylto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_8_5_5.C_ON=1'b0;
    defparam VSync_1_LC_8_5_5.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_8_5_5.LUT_INIT=16'b1111111111011111;
    LogicCell40 VSync_1_LC_8_5_5 (
            .in0(N__3969),
            .in1(N__3963),
            .in2(N__3909),
            .in3(N__3906),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5596),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_5_c_RNIB1PC_0_LC_8_5_6.C_ON=1'b0;
    defparam un5_visiblex_1_cry_5_c_RNIB1PC_0_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_5_c_RNIB1PC_0_LC_8_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_1_cry_5_c_RNIB1PC_0_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3822),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_6_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_6_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_6_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_LC_8_6_0 (
            .in0(_gnd_net_),
            .in1(N__3821),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05J52_LC_8_6_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05J52_LC_8_6_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05J52_LC_8_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05J52_LC_8_6_1 (
            .in0(_gnd_net_),
            .in1(N__4391),
            .in2(N__4239),
            .in3(N__3792),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4_c_RNI05JZ0Z52),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEO2_LC_8_6_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEO2_LC_8_6_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEO2_LC_8_6_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEO2_LC_8_6_2 (
            .in0(_gnd_net_),
            .in1(N__3789),
            .in2(N__3777),
            .in3(N__3768),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNIKUEOZ0Z2),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3NMD6_LC_8_6_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3NMD6_LC_8_6_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3NMD6_LC_8_6_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3NMD6_LC_8_6_3 (
            .in0(N__4733),
            .in1(N__4392),
            .in2(N__4383),
            .in3(N__4374),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_LC_8_6_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_LC_8_6_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_LC_8_6_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_LC_8_6_4 (
            .in0(_gnd_net_),
            .in1(N__4371),
            .in2(_gnd_net_),
            .in3(N__4365),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63),
            .ltout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUSZ0Z63_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_0_LC_8_6_5.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_0_LC_8_6_5.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_0_LC_8_6_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_7_c_RNIJUS63_0_LC_8_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4362),
            .in3(_gnd_net_),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIBKA_1_LC_8_6_6.C_ON=1'b0;
    defparam beamX_RNIBKA_1_LC_8_6_6.SEQ_MODE=4'b0000;
    defparam beamX_RNIBKA_1_LC_8_6_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_RNIBKA_1_LC_8_6_6 (
            .in0(N__4357),
            .in1(N__4308),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamX_RNIBKAZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_6_c_RNID4QC_0_LC_8_7_5.C_ON=1'b0;
    defparam un5_visiblex_1_cry_6_c_RNID4QC_0_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_6_c_RNID4QC_0_LC_8_7_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_1_cry_6_c_RNID4QC_0_LC_8_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4263),
            .lcout(un1_visiblex_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_1_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4847),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_1_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_9_1_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_9_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_9_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7H_LC_9_1_1 (
            .in0(_gnd_net_),
            .in1(N__4593),
            .in2(N__4639),
            .in3(N__4230),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_RNI0B7HZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFV81_LC_9_1_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFV81_LC_9_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFV81_LC_9_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFV81_LC_9_1_2 (
            .in0(_gnd_net_),
            .in1(N__4632),
            .in2(N__4227),
            .in3(N__4218),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3_c_RNINFVZ0Z81),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_9_1_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_9_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_9_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TK1_LC_9_1_3 (
            .in0(_gnd_net_),
            .in1(N__4707),
            .in2(N__4640),
            .in3(N__4701),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4_c_RNIH6TKZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI37VA3_LC_9_1_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI37VA3_LC_9_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI37VA3_LC_9_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_5_c_RNI37VA3_LC_9_1_4 (
            .in0(N__4913),
            .in1(N__4697),
            .in2(N__4686),
            .in3(N__4677),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_9_1_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_9_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_9_1_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_LC_9_1_5 (
            .in0(N__4674),
            .in1(N__4668),
            .in2(N__4641),
            .in3(N__4617),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVFZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_9_1_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_9_1_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_9_1_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_cry_6_c_RNIISVF_0_LC_9_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4614),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_1_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_1_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un40_sum_sbtinv_LC_9_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4610),
            .lcout(un1_beamY_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_fast_6_LC_9_2_2.C_ON=1'b0;
    defparam beamY_fast_6_LC_9_2_2.SEQ_MODE=4'b1000;
    defparam beamY_fast_6_LC_9_2_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 beamY_fast_6_LC_9_2_2 (
            .in0(N__4572),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamY_fastZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5600),
            .ce(N__4475),
            .sr(_gnd_net_));
    defparam beamY_6_LC_9_2_3.C_ON=1'b0;
    defparam beamY_6_LC_9_2_3.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_9_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_6_LC_9_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4571),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5600),
            .ce(N__4475),
            .sr(_gnd_net_));
    defparam beamY_2_LC_9_2_7.C_ON=1'b0;
    defparam beamY_2_LC_9_2_7.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_9_2_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_2_LC_9_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4508),
            .lcout(beamYZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5600),
            .ce(N__4475),
            .sr(_gnd_net_));
    defparam beamY_fast_2_LC_9_3_6.C_ON=1'b0;
    defparam beamY_fast_2_LC_9_3_6.SEQ_MODE=4'b1000;
    defparam beamY_fast_2_LC_9_3_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 beamY_fast_2_LC_9_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4512),
            .lcout(beamY_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5599),
            .ce(N__4470),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_5_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_5_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_5_0 (
            .in0(_gnd_net_),
            .in1(N__5492),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOS04_LC_9_5_1.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOS04_LC_9_5_1.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOS04_LC_9_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOS04_LC_9_5_1 (
            .in0(_gnd_net_),
            .in1(N__4788),
            .in2(N__4782),
            .in3(N__4773),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4_c_RNIPOSZ0Z04),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNP5_LC_9_5_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNP5_LC_9_5_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNP5_LC_9_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNP5_LC_9_5_2 (
            .in0(_gnd_net_),
            .in1(N__4734),
            .in2(N__4770),
            .in3(N__4761),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5_c_RNIFUNPZ0Z5),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_12_LC_9_5_3.C_ON=1'b1;
    defparam Pixel_1_RNO_12_LC_9_5_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_12_LC_9_5_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 Pixel_1_RNO_12_LC_9_5_3 (
            .in0(N__5539),
            .in1(N__4716),
            .in2(N__4746),
            .in3(N__4758),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0R6_LC_9_5_4.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0R6_LC_9_5_4.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0R6_LC_9_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0R6_LC_9_5_4 (
            .in0(_gnd_net_),
            .in1(N__4755),
            .in2(_gnd_net_),
            .in3(N__4749),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_cry_7_c_RNI1M0RZ0Z6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBV5_LC_9_5_7.C_ON=1'b0;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBV5_LC_9_5_7.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBV5_LC_9_5_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBV5_LC_9_5_7 (
            .in0(N__4745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4732),
            .lcout(un1_visiblex_if_generate_plus_mult1_un61_sum_cry_5_c_RNI7TBVZ0Z5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_1_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_1_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_1_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_1_0 (
            .in0(_gnd_net_),
            .in1(N__5184),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_1_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_11_1_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_11_1_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_11_1_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQ_LC_11_1_1 (
            .in0(_gnd_net_),
            .in1(N__4921),
            .in2(N__4821),
            .in3(N__4710),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_RNI1FUQZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_11_1_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_11_1_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_11_1_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQA1_LC_11_1_2 (
            .in0(_gnd_net_),
            .in1(N__4938),
            .in2(N__4926),
            .in3(N__4929),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3_c_RNIFCQAZ0Z1),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJ22_LC_11_1_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJ22_LC_11_1_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJ22_LC_11_1_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJ22_LC_11_1_3 (
            .in0(_gnd_net_),
            .in1(N__4925),
            .in2(N__4902),
            .in3(N__4890),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4_c_RNI7JJZ0Z22),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI5U736_LC_11_1_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI5U736_LC_11_1_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI5U736_LC_11_1_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_5_c_RNI5U736_LC_11_1_4 (
            .in0(N__5021),
            .in1(N__4887),
            .in2(N__4878),
            .in3(N__4866),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_LC_11_1_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_LC_11_1_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_LC_11_1_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_LC_11_1_5 (
            .in0(_gnd_net_),
            .in1(N__4863),
            .in2(_gnd_net_),
            .in3(N__4854),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILKZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_1_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_1_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_1_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un47_sum_sbtinv_LC_11_1_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4851),
            .lcout(un1_beamY_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_2_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_2_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_2_0 (
            .in0(_gnd_net_),
            .in1(N__5230),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONF4_LC_11_2_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONF4_LC_11_2_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONF4_LC_11_2_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONF4_LC_11_2_1 (
            .in0(_gnd_net_),
            .in1(N__5016),
            .in2(N__5154),
            .in3(N__4812),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_RNIEONFZ0Z4),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEV4_LC_11_2_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEV4_LC_11_2_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEV4_LC_11_2_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEV4_LC_11_2_2 (
            .in0(_gnd_net_),
            .in1(N__4809),
            .in2(N__5022),
            .in3(N__4803),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3_c_RNIVEEVZ0Z4),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBF5_LC_11_2_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBF5_LC_11_2_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBF5_LC_11_2_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBF5_LC_11_2_3 (
            .in0(_gnd_net_),
            .in1(N__5020),
            .in2(N__4800),
            .in3(N__4791),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4_c_RNIEEBFZ0Z5),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIA9BQC_LC_11_2_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIA9BQC_LC_11_2_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIA9BQC_LC_11_2_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_5_c_RNIA9BQC_LC_11_2_4 (
            .in0(N__4971),
            .in1(N__5043),
            .in2(N__4998),
            .in3(N__5037),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_LC_11_2_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_LC_11_2_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_LC_11_2_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_LC_11_2_5 (
            .in0(_gnd_net_),
            .in1(N__5034),
            .in2(_gnd_net_),
            .in3(N__5028),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6),
            .ltout(un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5JZ0Z6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_0_LC_11_2_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_0_LC_11_2_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_0_LC_11_2_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_cry_6_c_RNI3I5J6_0_LC_11_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5025),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_0_LC_11_2_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_0_LC_11_2_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_0_LC_11_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3ILK3_0_LC_11_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5015),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_3_0.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_3_0.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_3_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_3_0 (
            .in0(_gnd_net_),
            .in1(N__5819),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQ6_LC_11_3_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQ6_LC_11_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQ6_LC_11_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQ6_LC_11_3_1 (
            .in0(_gnd_net_),
            .in1(N__4972),
            .in2(N__5193),
            .in3(N__4989),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2_c_RNIJNKQZ0Z6),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85B_LC_11_3_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85B_LC_11_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85B_LC_11_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85B_LC_11_3_2 (
            .in0(_gnd_net_),
            .in1(N__4986),
            .in2(N__4977),
            .in3(N__4980),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3_c_RNIJC85BZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LB_LC_11_3_3.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LB_LC_11_3_3.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LB_LC_11_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LB_LC_11_3_3 (
            .in0(_gnd_net_),
            .in1(N__4976),
            .in2(N__4956),
            .in3(N__4947),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4_c_RNI550LBZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNI4ON1P_LC_11_3_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNI4ON1P_LC_11_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNI4ON1P_LC_11_3_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_5_c_RNI4ON1P_LC_11_3_4 (
            .in0(N__5875),
            .in1(N__4944),
            .in2(N__5253),
            .in3(N__5244),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSC_LC_11_3_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSC_LC_11_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSC_LC_11_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSC_LC_11_3_5 (
            .in0(_gnd_net_),
            .in1(N__5241),
            .in2(_gnd_net_),
            .in3(N__5235),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_cry_6_c_RNIFHPSCZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_11_3_6.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_11_3_6.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_11_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un61_sum_sbtinv_LC_11_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5232),
            .lcout(un1_beamY_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_3_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_3_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_3_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un54_sum_sbtinv_LC_11_3_7 (
            .in0(N__5182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un1_beamY_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_7_LC_11_4_4.C_ON=1'b0;
    defparam Pixel_1_RNO_7_LC_11_4_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_7_LC_11_4_4.LUT_INIT=16'b0011000101110011;
    LogicCell40 Pixel_1_RNO_7_LC_11_4_4 (
            .in0(N__5145),
            .in1(N__5073),
            .in2(N__5112),
            .in3(N__5054),
            .lcout(),
            .ltout(un19lto10_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_2_LC_11_4_5.C_ON=1'b0;
    defparam Pixel_1_RNO_2_LC_11_4_5.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_2_LC_11_4_5.LUT_INIT=16'b1010000101010000;
    LogicCell40 Pixel_1_RNO_2_LC_11_4_5 (
            .in0(N__5055),
            .in1(N__5111),
            .in2(N__5115),
            .in3(N__5502),
            .lcout(un19_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_11_5_0.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_11_5_0.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_11_5_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4_c_LC_11_5_0 (
            .in0(_gnd_net_),
            .in1(N__5107),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_13_LC_11_5_1.C_ON=1'b1;
    defparam Pixel_1_RNO_13_LC_11_5_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_13_LC_11_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_13_LC_11_5_1 (
            .in0(_gnd_net_),
            .in1(N__5522),
            .in2(N__5469),
            .in3(N__5067),
            .lcout(Pixel_1_RNOZ0Z_13),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVA_LC_11_5_2.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVA_LC_11_5_2.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVA_LC_11_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVA_LC_11_5_2 (
            .in0(_gnd_net_),
            .in1(N__5064),
            .in2(N__5544),
            .in3(N__5046),
            .lcout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5_c_RNIKICVAZ0),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_11_5_3.C_ON=1'b1;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_11_5_3.SEQ_MODE=4'b0000;
    defparam un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_11_5_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_11_5_3 (
            .in0(_gnd_net_),
            .in1(N__5523),
            .in2(N__5556),
            .in3(N__5540),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(un1_visiblex_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_6_LC_11_5_4.C_ON=1'b0;
    defparam Pixel_1_RNO_6_LC_11_5_4.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_6_LC_11_5_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 Pixel_1_RNO_6_LC_11_5_4 (
            .in0(_gnd_net_),
            .in1(N__5514),
            .in2(_gnd_net_),
            .in3(N__5505),
            .lcout(Pixel_1_RNOZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_visiblex_1_cry_4_c_RNI9UNC_0_LC_11_5_6.C_ON=1'b0;
    defparam un5_visiblex_1_cry_4_c_RNI9UNC_0_LC_11_5_6.SEQ_MODE=4'b0000;
    defparam un5_visiblex_1_cry_4_c_RNI9UNC_0_LC_11_5_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_visiblex_1_cry_4_c_RNI9UNC_0_LC_11_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5496),
            .lcout(un1_visiblex_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_11_5_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_11_5_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_11_5_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_11_5_7 (
            .in0(N__5456),
            .in1(N__5767),
            .in2(_gnd_net_),
            .in3(N__5350),
            .lcout(beamY_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_14_LC_12_3_0.C_ON=1'b1;
    defparam Pixel_1_RNO_14_LC_12_3_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_14_LC_12_3_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 Pixel_1_RNO_14_LC_12_3_0 (
            .in0(_gnd_net_),
            .in1(N__5768),
            .in2(_gnd_net_),
            .in3(N__5738),
            .lcout(G_6_i_a4_0_0),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9D_LC_12_3_1.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9D_LC_12_3_1.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9D_LC_12_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9D_LC_12_3_1 (
            .in0(_gnd_net_),
            .in1(N__5799),
            .in2(N__5876),
            .in3(N__5277),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_RNI4DJ9DZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00K_LC_12_3_2.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00K_LC_12_3_2.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00K_LC_12_3_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00K_LC_12_3_2 (
            .in0(_gnd_net_),
            .in1(N__5871),
            .in2(N__5274),
            .in3(N__5265),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3_c_RNI2K00KZ0),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_10_LC_12_3_3.C_ON=1'b1;
    defparam Pixel_1_RNO_10_LC_12_3_3.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_10_LC_12_3_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_1_RNO_10_LC_12_3_3 (
            .in0(_gnd_net_),
            .in1(N__5262),
            .in2(N__5877),
            .in3(N__5256),
            .lcout(Pixel_1_RNOZ0Z_10),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_12_3_4.C_ON=1'b1;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_12_3_4.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_12_3_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_12_3_4 (
            .in0(_gnd_net_),
            .in1(N__5883),
            .in2(N__5850),
            .in3(N__5867),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(un1_beamY_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAP_LC_12_3_5.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAP_LC_12_3_5.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAP_LC_12_3_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAP_LC_12_3_5 (
            .in0(_gnd_net_),
            .in1(N__5841),
            .in2(_gnd_net_),
            .in3(N__5835),
            .lcout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0),
            .ltout(un1_beamY_if_generate_plus_mult1_un75_sum_cry_6_c_RNI79DAPZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_9_LC_12_3_6.C_ON=1'b0;
    defparam Pixel_1_RNO_9_LC_12_3_6.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_9_LC_12_3_6.LUT_INIT=16'b0000100000000000;
    LogicCell40 Pixel_1_RNO_9_LC_12_3_6 (
            .in0(N__5832),
            .in1(N__5793),
            .in2(N__5826),
            .in3(N__5781),
            .lcout(N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_12_3_7.C_ON=1'b0;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_12_3_7.SEQ_MODE=4'b0000;
    defparam un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_12_3_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un1_beamY_if_generate_plus_mult1_un68_sum_sbtinv_LC_12_3_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5823),
            .lcout(un1_beamY_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_8_LC_12_4_0.C_ON=1'b0;
    defparam Pixel_1_RNO_8_LC_12_4_0.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_8_LC_12_4_0.LUT_INIT=16'b1110111111111111;
    LogicCell40 Pixel_1_RNO_8_LC_12_4_0 (
            .in0(N__5792),
            .in1(N__5780),
            .in2(N__5769),
            .in3(N__5745),
            .lcout(),
            .ltout(N_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_RNO_3_LC_12_4_1.C_ON=1'b0;
    defparam Pixel_1_RNO_3_LC_12_4_1.SEQ_MODE=4'b0000;
    defparam Pixel_1_RNO_3_LC_12_4_1.LUT_INIT=16'b0000000000110100;
    LogicCell40 Pixel_1_RNO_3_LC_12_4_1 (
            .in0(N__5739),
            .in1(N__5670),
            .in2(N__5664),
            .in3(N__5661),
            .lcout(),
            .ltout(un20_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_1_LC_12_4_2.C_ON=1'b0;
    defparam Pixel_1_LC_12_4_2.SEQ_MODE=4'b1000;
    defparam Pixel_1_LC_12_4_2.LUT_INIT=16'b0101101011001100;
    LogicCell40 Pixel_1_LC_12_4_2 (
            .in0(N__5655),
            .in1(N__5649),
            .in2(N__5637),
            .in3(N__5634),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5601),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
