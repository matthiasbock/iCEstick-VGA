// ******************************************************************************

// iCEcube Netlister

// Version:            2014.12.27052

// Build Date:         Dec  8 2014 15:16:04

// File Generated:     Jun 23 2015 21:37:58

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SimpleVGA" view "INTERFACE"

module SimpleVGA (
    VSyncDebug,
    PixelDebug,
    HSyncDebug,
    Clock12MHz,
    VSync,
    Pixel,
    HSync);

    output VSyncDebug;
    output PixelDebug;
    output HSyncDebug;
    input Clock12MHz;
    output VSync;
    output Pixel;
    output HSync;

    wire N__7874;
    wire N__7873;
    wire N__7872;
    wire N__7865;
    wire N__7864;
    wire N__7863;
    wire N__7856;
    wire N__7855;
    wire N__7854;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7838;
    wire N__7837;
    wire N__7836;
    wire N__7829;
    wire N__7828;
    wire N__7827;
    wire N__7820;
    wire N__7819;
    wire N__7818;
    wire N__7801;
    wire N__7800;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7782;
    wire N__7781;
    wire N__7780;
    wire N__7779;
    wire N__7778;
    wire N__7775;
    wire N__7774;
    wire N__7771;
    wire N__7770;
    wire N__7769;
    wire N__7768;
    wire N__7767;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7752;
    wire N__7749;
    wire N__7744;
    wire N__7741;
    wire N__7740;
    wire N__7737;
    wire N__7736;
    wire N__7735;
    wire N__7732;
    wire N__7731;
    wire N__7728;
    wire N__7727;
    wire N__7724;
    wire N__7723;
    wire N__7720;
    wire N__7715;
    wire N__7710;
    wire N__7707;
    wire N__7706;
    wire N__7705;
    wire N__7704;
    wire N__7703;
    wire N__7702;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7686;
    wire N__7671;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7625;
    wire N__7620;
    wire N__7615;
    wire N__7612;
    wire N__7607;
    wire N__7598;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7578;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7566;
    wire N__7561;
    wire N__7558;
    wire N__7555;
    wire N__7554;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7533;
    wire N__7530;
    wire N__7527;
    wire N__7522;
    wire N__7521;
    wire N__7520;
    wire N__7513;
    wire N__7510;
    wire N__7509;
    wire N__7508;
    wire N__7501;
    wire N__7498;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7488;
    wire N__7485;
    wire N__7482;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7467;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7459;
    wire N__7458;
    wire N__7457;
    wire N__7456;
    wire N__7455;
    wire N__7454;
    wire N__7451;
    wire N__7450;
    wire N__7449;
    wire N__7444;
    wire N__7441;
    wire N__7440;
    wire N__7439;
    wire N__7438;
    wire N__7437;
    wire N__7436;
    wire N__7435;
    wire N__7434;
    wire N__7423;
    wire N__7420;
    wire N__7415;
    wire N__7410;
    wire N__7405;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7375;
    wire N__7374;
    wire N__7373;
    wire N__7372;
    wire N__7371;
    wire N__7370;
    wire N__7369;
    wire N__7368;
    wire N__7367;
    wire N__7366;
    wire N__7365;
    wire N__7364;
    wire N__7363;
    wire N__7362;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7357;
    wire N__7356;
    wire N__7355;
    wire N__7354;
    wire N__7353;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7299;
    wire N__7298;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7294;
    wire N__7293;
    wire N__7292;
    wire N__7291;
    wire N__7290;
    wire N__7289;
    wire N__7288;
    wire N__7287;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7219;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7206;
    wire N__7205;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7167;
    wire N__7166;
    wire N__7165;
    wire N__7162;
    wire N__7159;
    wire N__7154;
    wire N__7147;
    wire N__7144;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7138;
    wire N__7137;
    wire N__7136;
    wire N__7135;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7119;
    wire N__7116;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7083;
    wire N__7080;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7062;
    wire N__7059;
    wire N__7056;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7020;
    wire N__7017;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7005;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6970;
    wire N__6969;
    wire N__6966;
    wire N__6965;
    wire N__6962;
    wire N__6957;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6927;
    wire N__6926;
    wire N__6923;
    wire N__6918;
    wire N__6913;
    wire N__6912;
    wire N__6907;
    wire N__6904;
    wire N__6903;
    wire N__6900;
    wire N__6897;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6853;
    wire N__6850;
    wire N__6849;
    wire N__6846;
    wire N__6845;
    wire N__6842;
    wire N__6837;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6807;
    wire N__6804;
    wire N__6803;
    wire N__6802;
    wire N__6801;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6785;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6771;
    wire N__6768;
    wire N__6765;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6751;
    wire N__6748;
    wire N__6747;
    wire N__6746;
    wire N__6745;
    wire N__6744;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6732;
    wire N__6727;
    wire N__6724;
    wire N__6715;
    wire N__6714;
    wire N__6713;
    wire N__6712;
    wire N__6711;
    wire N__6710;
    wire N__6707;
    wire N__6702;
    wire N__6697;
    wire N__6694;
    wire N__6685;
    wire N__6684;
    wire N__6683;
    wire N__6680;
    wire N__6679;
    wire N__6678;
    wire N__6675;
    wire N__6674;
    wire N__6671;
    wire N__6666;
    wire N__6661;
    wire N__6658;
    wire N__6649;
    wire N__6648;
    wire N__6647;
    wire N__6646;
    wire N__6643;
    wire N__6642;
    wire N__6639;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6619;
    wire N__6618;
    wire N__6617;
    wire N__6616;
    wire N__6611;
    wire N__6610;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6562;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6544;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6504;
    wire N__6503;
    wire N__6500;
    wire N__6495;
    wire N__6492;
    wire N__6489;
    wire N__6484;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6478;
    wire N__6477;
    wire N__6476;
    wire N__6475;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6460;
    wire N__6453;
    wire N__6442;
    wire N__6441;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6408;
    wire N__6405;
    wire N__6402;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6387;
    wire N__6386;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6367;
    wire N__6364;
    wire N__6361;
    wire N__6358;
    wire N__6355;
    wire N__6352;
    wire N__6349;
    wire N__6346;
    wire N__6345;
    wire N__6344;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6322;
    wire N__6319;
    wire N__6318;
    wire N__6315;
    wire N__6314;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6292;
    wire N__6289;
    wire N__6288;
    wire N__6285;
    wire N__6284;
    wire N__6283;
    wire N__6282;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6264;
    wire N__6253;
    wire N__6250;
    wire N__6249;
    wire N__6248;
    wire N__6245;
    wire N__6240;
    wire N__6239;
    wire N__6236;
    wire N__6235;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6220;
    wire N__6217;
    wire N__6212;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6171;
    wire N__6168;
    wire N__6165;
    wire N__6162;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6148;
    wire N__6145;
    wire N__6142;
    wire N__6141;
    wire N__6138;
    wire N__6135;
    wire N__6134;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6122;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6106;
    wire N__6103;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6071;
    wire N__6070;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6033;
    wire N__6030;
    wire N__6029;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6021;
    wire N__6018;
    wire N__6011;
    wire N__6004;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5992;
    wire N__5989;
    wire N__5988;
    wire N__5985;
    wire N__5984;
    wire N__5981;
    wire N__5976;
    wire N__5971;
    wire N__5970;
    wire N__5969;
    wire N__5966;
    wire N__5961;
    wire N__5956;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5898;
    wire N__5897;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5885;
    wire N__5882;
    wire N__5875;
    wire N__5872;
    wire N__5871;
    wire N__5868;
    wire N__5867;
    wire N__5862;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5852;
    wire N__5845;
    wire N__5842;
    wire N__5841;
    wire N__5840;
    wire N__5837;
    wire N__5832;
    wire N__5827;
    wire N__5824;
    wire N__5823;
    wire N__5818;
    wire N__5815;
    wire N__5812;
    wire N__5809;
    wire N__5808;
    wire N__5807;
    wire N__5806;
    wire N__5803;
    wire N__5798;
    wire N__5795;
    wire N__5792;
    wire N__5789;
    wire N__5782;
    wire N__5781;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5745;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5679;
    wire N__5678;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5656;
    wire N__5655;
    wire N__5654;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5641;
    wire N__5632;
    wire N__5629;
    wire N__5628;
    wire N__5627;
    wire N__5624;
    wire N__5623;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5611;
    wire N__5608;
    wire N__5599;
    wire N__5598;
    wire N__5597;
    wire N__5596;
    wire N__5595;
    wire N__5592;
    wire N__5589;
    wire N__5584;
    wire N__5581;
    wire N__5572;
    wire N__5569;
    wire N__5568;
    wire N__5567;
    wire N__5566;
    wire N__5565;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5550;
    wire N__5547;
    wire N__5536;
    wire N__5535;
    wire N__5534;
    wire N__5533;
    wire N__5532;
    wire N__5529;
    wire N__5528;
    wire N__5527;
    wire N__5526;
    wire N__5523;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5507;
    wire N__5504;
    wire N__5491;
    wire N__5490;
    wire N__5489;
    wire N__5488;
    wire N__5487;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5472;
    wire N__5469;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5448;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5442;
    wire N__5441;
    wire N__5438;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5370;
    wire N__5365;
    wire N__5364;
    wire N__5363;
    wire N__5362;
    wire N__5361;
    wire N__5358;
    wire N__5355;
    wire N__5352;
    wire N__5347;
    wire N__5338;
    wire N__5337;
    wire N__5336;
    wire N__5335;
    wire N__5332;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5295;
    wire N__5294;
    wire N__5293;
    wire N__5292;
    wire N__5289;
    wire N__5284;
    wire N__5279;
    wire N__5272;
    wire N__5271;
    wire N__5268;
    wire N__5265;
    wire N__5262;
    wire N__5257;
    wire N__5256;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5208;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5190;
    wire N__5189;
    wire N__5186;
    wire N__5185;
    wire N__5182;
    wire N__5175;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5151;
    wire N__5150;
    wire N__5145;
    wire N__5142;
    wire N__5139;
    wire N__5136;
    wire N__5133;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5118;
    wire N__5115;
    wire N__5114;
    wire N__5111;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5089;
    wire N__5088;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5070;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5028;
    wire N__5027;
    wire N__5024;
    wire N__5023;
    wire N__5022;
    wire N__5019;
    wire N__5016;
    wire N__5007;
    wire N__5002;
    wire N__4999;
    wire N__4996;
    wire N__4995;
    wire N__4990;
    wire N__4989;
    wire N__4986;
    wire N__4983;
    wire N__4980;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4963;
    wire N__4960;
    wire N__4957;
    wire N__4956;
    wire N__4951;
    wire N__4948;
    wire N__4945;
    wire N__4942;
    wire N__4941;
    wire N__4938;
    wire N__4935;
    wire N__4930;
    wire N__4927;
    wire N__4924;
    wire N__4921;
    wire N__4918;
    wire N__4915;
    wire N__4912;
    wire N__4909;
    wire N__4906;
    wire N__4903;
    wire N__4900;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4888;
    wire N__4887;
    wire N__4884;
    wire N__4883;
    wire N__4882;
    wire N__4875;
    wire N__4872;
    wire N__4867;
    wire N__4864;
    wire N__4861;
    wire N__4858;
    wire N__4855;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4840;
    wire N__4837;
    wire N__4834;
    wire N__4831;
    wire N__4828;
    wire N__4825;
    wire N__4822;
    wire N__4819;
    wire N__4816;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4804;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4794;
    wire N__4791;
    wire N__4790;
    wire N__4787;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4775;
    wire N__4768;
    wire N__4765;
    wire N__4762;
    wire N__4759;
    wire N__4756;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4729;
    wire N__4726;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4698;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4672;
    wire N__4669;
    wire N__4666;
    wire N__4663;
    wire N__4660;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4647;
    wire N__4644;
    wire N__4641;
    wire N__4636;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4608;
    wire N__4605;
    wire N__4604;
    wire N__4603;
    wire N__4596;
    wire N__4593;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4552;
    wire N__4549;
    wire N__4546;
    wire N__4543;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4533;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4500;
    wire N__4495;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4459;
    wire N__4456;
    wire N__4453;
    wire N__4450;
    wire N__4447;
    wire N__4444;
    wire N__4441;
    wire N__4438;
    wire N__4435;
    wire N__4432;
    wire N__4431;
    wire N__4428;
    wire N__4427;
    wire N__4426;
    wire N__4419;
    wire N__4416;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4399;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4387;
    wire N__4384;
    wire N__4381;
    wire N__4378;
    wire N__4377;
    wire N__4376;
    wire N__4375;
    wire N__4372;
    wire N__4365;
    wire N__4362;
    wire N__4359;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4344;
    wire N__4343;
    wire N__4342;
    wire N__4339;
    wire N__4336;
    wire N__4333;
    wire N__4330;
    wire N__4321;
    wire N__4318;
    wire N__4315;
    wire N__4312;
    wire N__4311;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4300;
    wire N__4299;
    wire N__4296;
    wire N__4287;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4242;
    wire N__4239;
    wire N__4238;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4225;
    wire N__4216;
    wire N__4213;
    wire N__4212;
    wire N__4211;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4198;
    wire N__4189;
    wire N__4188;
    wire N__4187;
    wire N__4182;
    wire N__4179;
    wire N__4176;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4155;
    wire N__4154;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4141;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4123;
    wire N__4122;
    wire N__4121;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4105;
    wire N__4102;
    wire N__4099;
    wire N__4096;
    wire N__4093;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4039;
    wire N__4038;
    wire N__4035;
    wire N__4032;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4015;
    wire N__4012;
    wire N__4009;
    wire N__4008;
    wire N__4007;
    wire N__4004;
    wire N__3999;
    wire N__3994;
    wire N__3991;
    wire N__3990;
    wire N__3989;
    wire N__3986;
    wire N__3981;
    wire N__3976;
    wire N__3973;
    wire N__3970;
    wire N__3967;
    wire N__3964;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3952;
    wire N__3949;
    wire N__3948;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3936;
    wire N__3933;
    wire N__3930;
    wire N__3927;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3879;
    wire N__3878;
    wire N__3875;
    wire N__3874;
    wire N__3865;
    wire N__3862;
    wire N__3859;
    wire N__3856;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3846;
    wire N__3843;
    wire N__3840;
    wire N__3835;
    wire N__3832;
    wire N__3829;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3808;
    wire N__3805;
    wire N__3802;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3784;
    wire N__3781;
    wire N__3778;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3730;
    wire N__3727;
    wire N__3724;
    wire N__3721;
    wire N__3718;
    wire N__3715;
    wire N__3712;
    wire N__3709;
    wire N__3706;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire \Clock50MHz.PixelClock ;
    wire Clock12MHz_c;
    wire VCCG0;
    wire bfn_4_3_0_;
    wire r_if_generate_plus_mult1_un68_sum_cry_2;
    wire r_if_generate_plus_mult1_un68_sum_cry_3;
    wire r_if_generate_plus_mult1_un68_sum_cry_4;
    wire r_if_generate_plus_mult1_un61_sum_i_5;
    wire r_if_generate_plus_mult1_un61_sum_i_0;
    wire bfn_4_5_0_;
    wire if_generate_plus_mult1_un61_sum_cry_3_s_0;
    wire r_if_generate_plus_mult1_un61_sum_cry_2;
    wire r_if_generate_plus_mult1_un68_sum_axbZ0Z_5;
    wire r_if_generate_plus_mult1_un61_sum_cry_3;
    wire r_if_generate_plus_mult1_un61_sum_cry_4;
    wire bfn_4_6_0_;
    wire if_generate_plus_mult1_un54_sum_cry_3_s_0;
    wire r_if_generate_plus_mult1_un54_sum_cry_2;
    wire r_if_generate_plus_mult1_un61_sum_axbZ0Z_5;
    wire r_if_generate_plus_mult1_un54_sum_cry_3;
    wire r_if_generate_plus_mult1_un54_sum_cry_4;
    wire bfn_4_7_0_;
    wire if_generate_plus_mult1_un47_sum_cry_3_s;
    wire r_if_generate_plus_mult1_un47_sum_cry_2;
    wire r_if_generate_plus_mult1_un54_sum_axbZ0Z_5;
    wire r_if_generate_plus_mult1_un47_sum_cry_3;
    wire r_if_generate_plus_mult1_un47_sum_cry_4;
    wire visibleYZ0Z_6;
    wire bfn_4_9_0_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1_cascade_;
    wire visibleYZ0Z_7;
    wire bfn_4_10_0_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450QZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9MZ0Z01;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDOZ0Z01;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0_cascade_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_7;
    wire visibleY_RNINQ3DZ0Z_8;
    wire bfn_5_2_0_;
    wire G_251;
    wire r_if_generate_plus_mult1_un82_sum_cry_2;
    wire G_252;
    wire r_if_generate_plus_mult1_un82_sum_cry_3;
    wire r_if_generate_plus_mult1_un82_sum_cry_4;
    wire G_250;
    wire bfn_5_3_0_;
    wire r_if_generate_plus_mult1_un68_sum_i_0;
    wire if_generate_plus_mult1_un75_sum_cry_3_s;
    wire r_if_generate_plus_mult1_un75_sum_cry_2;
    wire r_if_generate_plus_mult1_un68_sum_i_5;
    wire if_generate_plus_mult1_un68_sum_cry_3_s_0;
    wire r_if_generate_plus_mult1_un82_sum_axbZ0Z_5;
    wire r_if_generate_plus_mult1_un75_sum_cry_3;
    wire r_if_generate_plus_mult1_un75_sum_axbZ0Z_5;
    wire r_if_generate_plus_mult1_un75_sum_cry_4;
    wire bfn_5_4_0_;
    wire r_if_generate_plus_mult1_un75_sum;
    wire un5_vy_cry_0;
    wire r_if_generate_plus_mult1_un68_sum;
    wire un5_vy_cry_1;
    wire r_if_generate_plus_mult1_un61_sum;
    wire un5_vy_cry_2;
    wire un5_vy_cry_3;
    wire un5_vy_cry_4;
    wire un5_vy_cry_5;
    wire un5_vy_cry_6;
    wire if_generate_plus_mult1_un61_sum_s_5;
    wire if_generate_plus_mult1_un68_sum_s_5;
    wire r_if_generate_plus_mult1_un54_sum;
    wire r_if_generate_plus_mult1_un54_sum_i_0;
    wire r_if_generate_plus_mult1_un54_sum_i_5;
    wire if_generate_plus_mult1_un54_sum_s_5_0;
    wire un7_r_1;
    wire r_if_generate_plus_mult1_un47_sum;
    wire r_if_generate_plus_mult1_un47_sum_i_0;
    wire un5_vy_cry_6_c_RNIG9KKZ0;
    wire if_generate_plus_mult1_un47_sum_axb_4_l_ofx;
    wire un5_vy_cry_6_c_RNI9MAAZ0;
    wire N_7_i;
    wire if_generate_plus_mult1_un47_sum_s_5;
    wire r_if_generate_plus_mult1_un47_sum_i_5;
    wire un5_vy_cry_5_c_RNI7J9AZ0;
    wire un5_vy_i_24;
    wire bfn_5_8_0_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0_cascade_;
    wire visibleYZ0Z_4;
    wire visibleYZ0Z_5;
    wire bfn_5_9_0_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_i_0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSVZ0Z1;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71EZ0Z1;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0VZ0Z33;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5TZ0Z1;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4JZ0Z3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5KZ0Z3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_axb_7;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_axb_7;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3_cascade_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_7;
    wire visibleYZ0Z_8;
    wire bfn_5_10_0_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6;
    wire visibleYZ0Z_9;
    wire visibleY_RNIOR3DZ0Z_9;
    wire bfn_5_11_0_;
    wire c_if_generate_plus_mult1_un61_sum_iZ0;
    wire c_if_generate_plus_mult1_un68_sum_cry_1;
    wire c_if_generate_plus_mult1_un68_sum_cry_2;
    wire c_if_generate_plus_mult1_un68_sum_cry_3;
    wire c_if_generate_plus_mult1_un68_sum_cry_4;
    wire bfn_5_12_0_;
    wire if_generate_plus_mult1_un61_sum_cry_2_s;
    wire c_if_generate_plus_mult1_un61_sum_cry_1;
    wire if_generate_plus_mult1_un61_sum_cry_3_s;
    wire c_if_generate_plus_mult1_un61_sum_cry_2;
    wire c_if_generate_plus_mult1_un68_sum_axbZ0Z_5;
    wire c_if_generate_plus_mult1_un61_sum_cry_3;
    wire c_if_generate_plus_mult1_un61_sum_cry_4;
    wire bfn_6_3_0_;
    wire un21_beamy_cry_1;
    wire un21_beamy_cry_1_THRU_CRY_0_THRU_CO;
    wire un21_beamy_cry_1_THRU_CRY_1_THRU_CO;
    wire un21_beamy_cry_1_THRU_CRY_2_THRU_CO;
    wire un21_beamy_cry_1_THRU_CRY_3_THRU_CO;
    wire un21_beamy_cry_1_THRU_CRY_4_THRU_CO;
    wire GNDG0;
    wire un21_beamy_cry_1_THRU_CRY_5_THRU_CO;
    wire un21_beamy_cry_1_THRU_CRY_6_THRU_CO;
    wire bfn_6_4_0_;
    wire un21_beamy_cry_2;
    wire un21_beamy_cry_3;
    wire un21_beamy_cry_4;
    wire un21_beamy_cry_5;
    wire un21_beamy_cry_6;
    wire un21_beamy_cry_7;
    wire un21_beamy_cry_8;
    wire if_generate_plus_mult1_un82_sum_s_5;
    wire un7_r_4;
    wire if_generate_plus_mult1_un75_sum_s_5;
    wire bfn_6_7_0_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_7;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41_cascade_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7CZ0Z11;
    wire Pixel_RNOZ0Z_7;
    wire visibleYZ0Z_3;
    wire bfn_6_8_0_;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000BZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73PZ0Z94;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SEZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQZ0Z56;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OGZ0;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUTZ0Z97;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_7;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_axb_7;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_axb_7;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0;
    wire bfn_6_9_0_;
    wire un5_vx_cry_0;
    wire un5_vx_cry_1;
    wire un5_vx_cry_2;
    wire c_if_generate_plus_mult1_un61_sum;
    wire un5_vx_cry_3;
    wire un5_vx_cry_4;
    wire un5_vx_cry_5;
    wire un5_vx_cry_6;
    wire un5_vx_cry_7;
    wire bfn_6_10_0_;
    wire un5_vx_cry_8;
    wire CO3_0_cascade_;
    wire N_14;
    wire N_3_0_cascade_;
    wire c_if_generate_plus_mult1_un75_sum;
    wire bfn_6_11_0_;
    wire c_if_generate_plus_mult1_un75_sum_cry_1;
    wire if_generate_plus_mult1_un68_sum_cry_2_s;
    wire c_if_generate_plus_mult1_un75_sum_cry_2;
    wire G_253;
    wire if_generate_plus_mult1_un68_sum_cry_3_s;
    wire c_if_generate_plus_mult1_un75_sum_cry_3;
    wire un9_r_0lto2;
    wire c_if_generate_plus_mult1_un75_sum_axbZ0Z_5;
    wire c_if_generate_plus_mult1_un75_sum_cry_4;
    wire un9_r_1lt6_0;
    wire c_if_generate_plus_mult1_un68_sum;
    wire c_if_generate_plus_mult1_un68_sum_iZ0;
    wire un9_r_0lto3;
    wire un9_r_0lto3_i;
    wire N_404_i;
    wire c_if_generate_plus_mult1_un54_sum_i_5;
    wire beamY_RNI9DLCZ0Z_2;
    wire beamYZ0Z_0;
    wire un5_beamx_5;
    wire un1_beamy_4_cascade_;
    wire un5_beamx_3;
    wire beamYZ0Z_1;
    wire un1_beamy_4;
    wire un8_beamy_2;
    wire un1_beamylto9_2_cascade_;
    wire VSync_c;
    wire beamYZ0Z_6;
    wire beamYZ0Z_5;
    wire un4_beamylt6_cascade_;
    wire beamYZ0Z_9;
    wire beamYZ0Z_8;
    wire un4_beamylt8_0_cascade_;
    wire beamYZ0Z_7;
    wire un5_vy;
    wire beamYZ0Z_4;
    wire un8_beamylto9_1;
    wire beamYZ0Z_3;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41;
    wire Pixel_RNOZ0Z_5_cascade_;
    wire N_45_cascade_;
    wire N_76;
    wire TextOutputEnabledZ0;
    wire N_74_i_cascade_;
    wire Pixel_c;
    wire INVPixelZ0C_net;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0;
    wire visibleYZ0Z_1;
    wire visibleYZ0Z_2;
    wire chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0;
    wire Pixel_RNOZ0Z_6;
    wire un13_beamylt7_cascade_;
    wire OutputEnabledZ0;
    wire un18_beamylt4;
    wire un18_beamylto9_2_cascade_;
    wire un8_beamy;
    wire un18_beamylt10_0_cascade_;
    wire un4_beamy_0;
    wire un15_beamy_2;
    wire un13_beamylt7;
    wire un15_beamy_2_cascade_;
    wire beamX_RNISO4TZ0Z_7;
    wire bfn_7_8_0_;
    wire un8_beamx_cry_1;
    wire un8_beamx_cry_2;
    wire un8_beamx_cry_3;
    wire un8_beamx_cry_4;
    wire un8_beamx_cry_5;
    wire un8_beamx_cry_6;
    wire beamXZ0Z_8;
    wire un8_beamx_cry_7;
    wire un8_beamx_cry_8;
    wire beamXZ0Z_9;
    wire bfn_7_9_0_;
    wire un8_beamx_cry_9;
    wire un5_vx_i_25_cascade_;
    wire bfn_7_10_0_;
    wire un5_vx_i_0_25;
    wire c_if_generate_plus_mult1_un47_sum_1_cry_1;
    wire c_if_generate_plus_mult1_un47_sum_0_axb_5_i;
    wire N_13_0_i;
    wire c_if_generate_plus_mult1_un47_sum_1_cry_2;
    wire if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx;
    wire c_if_generate_plus_mult1_un47_sum_1_cry_3;
    wire c_if_generate_plus_mult1_un47_sum_1_cry_4;
    wire c_if_generate_plus_mult1_un47_sum_0_0;
    wire c_if_generate_plus_mult1_un47_sum1_4;
    wire N_18_cascade_;
    wire c_if_generate_plus_mult1_un47_sum1_3;
    wire c_if_generate_plus_mult1_un47_sum1_5;
    wire c_if_generate_plus_mult1_un47_sum1_0;
    wire bfn_7_12_0_;
    wire if_generate_plus_mult1_un54_sum_axb_2_l_fx;
    wire if_generate_plus_mult1_un54_sum_cry_2_s;
    wire c_if_generate_plus_mult1_un54_sum_cry_1;
    wire if_generate_plus_mult1_un54_sum_axb_3_l_fx;
    wire if_generate_plus_mult1_un47_sum_m_2;
    wire if_generate_plus_mult1_un54_sum_cry_3_s;
    wire c_if_generate_plus_mult1_un54_sum_cry_2;
    wire N_18;
    wire if_generate_plus_mult1_un54_sum_axb_4_l_fx;
    wire c_if_generate_plus_mult1_un61_sum_axbZ0Z_5;
    wire c_if_generate_plus_mult1_un54_sum_cry_3;
    wire c_if_generate_plus_mult1_un54_sum_axbZ0Z_5;
    wire c_if_generate_plus_mult1_un54_sum_cry_4;
    wire if_generate_plus_mult1_un54_sum_s_5;
    wire bfn_8_7_0_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i_8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_6;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7;
    wire N_84;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0_cascade_;
    wire N_53;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0;
    wire Pixel_RNOZ0Z_8;
    wire visibleXZ0Z_4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0;
    wire N_81;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i;
    wire beamXZ0Z_2;
    wire beamXZ0Z_1;
    wire un3_beamx_5_cascade_;
    wire un5_vx;
    wire un3_beamx_7_cascade_;
    wire beamX_RNI5457Z0Z_5;
    wire beamXZ0Z_6;
    wire beamXZ0Z_4;
    wire beamXZ0Z_5;
    wire beamXZ0Z_3;
    wire c_if_generate_plus_mult1_un47_sum_1;
    wire bfn_8_9_0_;
    wire if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx;
    wire un5_vx_i_25;
    wire c_if_generate_plus_mult1_un47_sum0_2;
    wire c_if_generate_plus_mult1_un47_sum_0_cry_1;
    wire if_generate_plus_mult1_un47_sum_0_cry_3_ma;
    wire if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx;
    wire c_if_generate_plus_mult1_un47_sum0_3;
    wire c_if_generate_plus_mult1_un47_sum_0_cry_2;
    wire N_186_0_i;
    wire c_if_generate_plus_mult1_un47_sum0_4;
    wire c_if_generate_plus_mult1_un47_sum_0_cry_3;
    wire c_if_generate_plus_mult1_un47_sum_0_cry_4;
    wire c_if_generate_plus_mult1_un47_sum0_5;
    wire un5_vx_cry_6_c_RNI59BZ0;
    wire bfn_8_10_0_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412_cascade_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i;
    wire N_3_0;
    wire if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx;
    wire visibleXZ0Z_8;
    wire bfn_8_11_0_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29RZ0Z21;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKVZ0;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_axb_8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i_8;
    wire visibleXZ0Z_5;
    wire bfn_9_8_0_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56BZ0Z05;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNICZ0Z7997;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_axb_8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEAZ0Z08;
    wire beamXZ0Z_10;
    wire un1_beamx_2;
    wire beamXZ0Z_7;
    wire un1_beamxlt10_0;
    wire HSync_c;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i;
    wire visibleXZ0Z_6;
    wire bfn_9_9_0_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTKZ0Z2;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BDZ0Z1;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19MZ0Z3;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i_8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMKZ0Z642;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_axb_8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_axb_8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4_cascade_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i_8;
    wire visibleXZ0Z_7;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i;
    wire CO3_0;
    wire PixelClock_g;
    wire un15_beamy_g;
    wire bfn_9_11_0_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8PZ0Z8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQZ0Z8;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7;
    wire visibleXZ0Z_9;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i;
    wire CONSTANT_ONE_NET;
    wire bfn_9_12_0_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0_cascade_;
    wire chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i_8;
    wire G_255_cascade_;
    wire G_256;
    wire CharacterDisplay__decfrac8;
    wire G_255;
    wire G_254;
    wire _gnd_net_;

    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \Clock50MHz.PLL_inst .TEST_MODE=1'b0;
    defparam \Clock50MHz.PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \Clock50MHz.PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \Clock50MHz.PLL_inst .FILTER_RANGE=3'b001;
    defparam \Clock50MHz.PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \Clock50MHz.PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \Clock50MHz.PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \Clock50MHz.PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \Clock50MHz.PLL_inst .DIVR=4'b0000;
    defparam \Clock50MHz.PLL_inst .DIVQ=3'b100;
    defparam \Clock50MHz.PLL_inst .DIVF=7'b1000010;
    defparam \Clock50MHz.PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \Clock50MHz.PLL_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\Clock50MHz.PixelClock ),
            .REFERENCECLK(N__3688),
            .RESETB(N__7752),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam PixelDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD PixelDebug_obuf_iopad (
            .OE(N__7874),
            .DIN(N__7873),
            .DOUT(N__7872),
            .PACKAGEPIN(PixelDebug));
    defparam PixelDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PixelDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PixelDebug_obuf_preio (
            .PADOEN(N__7874),
            .PADOUT(N__7873),
            .PADIN(N__7872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7533),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSync_obuf_iopad (
            .OE(N__7865),
            .DIN(N__7864),
            .DOUT(N__7863),
            .PACKAGEPIN(VSync));
    defparam VSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSync_obuf_preio (
            .PADOEN(N__7865),
            .PADOUT(N__7864),
            .PADIN(N__7863),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5238),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSync_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSync_obuf_iopad (
            .OE(N__7856),
            .DIN(N__7855),
            .DOUT(N__7854),
            .PACKAGEPIN(HSync));
    defparam HSync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSync_obuf_preio (
            .PADOEN(N__7856),
            .PADOUT(N__7855),
            .PADIN(N__7854),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7092),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Clock12MHz_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Clock12MHz_ibuf_iopad (
            .OE(N__7847),
            .DIN(N__7846),
            .DOUT(N__7845),
            .PACKAGEPIN(Clock12MHz));
    defparam Clock12MHz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam Clock12MHz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO Clock12MHz_ibuf_preio (
            .PADOEN(N__7847),
            .PADOUT(N__7846),
            .PADIN(N__7845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(Clock12MHz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam HSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD HSyncDebug_obuf_iopad (
            .OE(N__7838),
            .DIN(N__7837),
            .DOUT(N__7836),
            .PACKAGEPIN(HSyncDebug));
    defparam HSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HSyncDebug_obuf_preio (
            .PADOEN(N__7838),
            .PADOUT(N__7837),
            .PADIN(N__7836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7099),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam Pixel_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD Pixel_obuf_iopad (
            .OE(N__7829),
            .DIN(N__7828),
            .DOUT(N__7827),
            .PACKAGEPIN(Pixel));
    defparam Pixel_obuf_preio.NEG_TRIGGER=1'b0;
    defparam Pixel_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO Pixel_obuf_preio (
            .PADOEN(N__7829),
            .PADOUT(N__7828),
            .PADIN(N__7827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5386),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VSyncDebug_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD VSyncDebug_obuf_iopad (
            .OE(N__7820),
            .DIN(N__7819),
            .DOUT(N__7818),
            .PACKAGEPIN(VSyncDebug));
    defparam VSyncDebug_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VSyncDebug_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VSyncDebug_obuf_preio (
            .PADOEN(N__7820),
            .PADOUT(N__7819),
            .PADIN(N__7818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1699 (
            .O(N__7801),
            .I(N__7795));
    InMux I__1698 (
            .O(N__7800),
            .I(N__7795));
    LocalMux I__1697 (
            .O(N__7795),
            .I(visibleXZ0Z_9));
    CascadeMux I__1696 (
            .O(N__7792),
            .I(N__7789));
    InMux I__1695 (
            .O(N__7789),
            .I(N__7786));
    LocalMux I__1694 (
            .O(N__7786),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i));
    CascadeMux I__1693 (
            .O(N__7783),
            .I(N__7775));
    CascadeMux I__1692 (
            .O(N__7782),
            .I(N__7771));
    CascadeMux I__1691 (
            .O(N__7781),
            .I(N__7763));
    CascadeMux I__1690 (
            .O(N__7780),
            .I(N__7760));
    CascadeMux I__1689 (
            .O(N__7779),
            .I(N__7757));
    CascadeMux I__1688 (
            .O(N__7778),
            .I(N__7754));
    InMux I__1687 (
            .O(N__7775),
            .I(N__7749));
    InMux I__1686 (
            .O(N__7774),
            .I(N__7744));
    InMux I__1685 (
            .O(N__7771),
            .I(N__7744));
    InMux I__1684 (
            .O(N__7770),
            .I(N__7741));
    CascadeMux I__1683 (
            .O(N__7769),
            .I(N__7737));
    CascadeMux I__1682 (
            .O(N__7768),
            .I(N__7732));
    CascadeMux I__1681 (
            .O(N__7767),
            .I(N__7728));
    CascadeMux I__1680 (
            .O(N__7766),
            .I(N__7724));
    InMux I__1679 (
            .O(N__7763),
            .I(N__7720));
    InMux I__1678 (
            .O(N__7760),
            .I(N__7715));
    InMux I__1677 (
            .O(N__7757),
            .I(N__7715));
    InMux I__1676 (
            .O(N__7754),
            .I(N__7710));
    InMux I__1675 (
            .O(N__7753),
            .I(N__7710));
    IoInMux I__1674 (
            .O(N__7752),
            .I(N__7707));
    LocalMux I__1673 (
            .O(N__7749),
            .I(N__7697));
    LocalMux I__1672 (
            .O(N__7744),
            .I(N__7697));
    LocalMux I__1671 (
            .O(N__7741),
            .I(N__7694));
    InMux I__1670 (
            .O(N__7740),
            .I(N__7691));
    InMux I__1669 (
            .O(N__7737),
            .I(N__7686));
    InMux I__1668 (
            .O(N__7736),
            .I(N__7686));
    InMux I__1667 (
            .O(N__7735),
            .I(N__7671));
    InMux I__1666 (
            .O(N__7732),
            .I(N__7671));
    InMux I__1665 (
            .O(N__7731),
            .I(N__7671));
    InMux I__1664 (
            .O(N__7728),
            .I(N__7671));
    InMux I__1663 (
            .O(N__7727),
            .I(N__7671));
    InMux I__1662 (
            .O(N__7724),
            .I(N__7671));
    InMux I__1661 (
            .O(N__7723),
            .I(N__7671));
    LocalMux I__1660 (
            .O(N__7720),
            .I(N__7664));
    LocalMux I__1659 (
            .O(N__7715),
            .I(N__7664));
    LocalMux I__1658 (
            .O(N__7710),
            .I(N__7664));
    LocalMux I__1657 (
            .O(N__7707),
            .I(N__7661));
    InMux I__1656 (
            .O(N__7706),
            .I(N__7658));
    CascadeMux I__1655 (
            .O(N__7705),
            .I(N__7655));
    CascadeMux I__1654 (
            .O(N__7704),
            .I(N__7652));
    CascadeMux I__1653 (
            .O(N__7703),
            .I(N__7649));
    CascadeMux I__1652 (
            .O(N__7702),
            .I(N__7646));
    Span4Mux_v I__1651 (
            .O(N__7697),
            .I(N__7643));
    Span4Mux_v I__1650 (
            .O(N__7694),
            .I(N__7636));
    LocalMux I__1649 (
            .O(N__7691),
            .I(N__7636));
    LocalMux I__1648 (
            .O(N__7686),
            .I(N__7636));
    LocalMux I__1647 (
            .O(N__7671),
            .I(N__7633));
    Span4Mux_v I__1646 (
            .O(N__7664),
            .I(N__7630));
    IoSpan4Mux I__1645 (
            .O(N__7661),
            .I(N__7625));
    LocalMux I__1644 (
            .O(N__7658),
            .I(N__7625));
    InMux I__1643 (
            .O(N__7655),
            .I(N__7620));
    InMux I__1642 (
            .O(N__7652),
            .I(N__7620));
    InMux I__1641 (
            .O(N__7649),
            .I(N__7615));
    InMux I__1640 (
            .O(N__7646),
            .I(N__7615));
    Span4Mux_v I__1639 (
            .O(N__7643),
            .I(N__7612));
    Span4Mux_v I__1638 (
            .O(N__7636),
            .I(N__7607));
    Span4Mux_h I__1637 (
            .O(N__7633),
            .I(N__7607));
    Span4Mux_v I__1636 (
            .O(N__7630),
            .I(N__7598));
    Span4Mux_s3_v I__1635 (
            .O(N__7625),
            .I(N__7598));
    LocalMux I__1634 (
            .O(N__7620),
            .I(N__7598));
    LocalMux I__1633 (
            .O(N__7615),
            .I(N__7598));
    Odrv4 I__1632 (
            .O(N__7612),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1631 (
            .O(N__7607),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1630 (
            .O(N__7598),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1629 (
            .O(N__7591),
            .I(N__7588));
    InMux I__1628 (
            .O(N__7588),
            .I(N__7585));
    LocalMux I__1627 (
            .O(N__7585),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO));
    InMux I__1626 (
            .O(N__7582),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6));
    InMux I__1625 (
            .O(N__7579),
            .I(N__7573));
    InMux I__1624 (
            .O(N__7578),
            .I(N__7573));
    LocalMux I__1623 (
            .O(N__7573),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0));
    CascadeMux I__1622 (
            .O(N__7570),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0_cascade_));
    InMux I__1621 (
            .O(N__7567),
            .I(N__7561));
    InMux I__1620 (
            .O(N__7566),
            .I(N__7561));
    LocalMux I__1619 (
            .O(N__7561),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i_8));
    CascadeMux I__1618 (
            .O(N__7558),
            .I(G_255_cascade_));
    InMux I__1617 (
            .O(N__7555),
            .I(N__7549));
    InMux I__1616 (
            .O(N__7554),
            .I(N__7549));
    LocalMux I__1615 (
            .O(N__7549),
            .I(G_256));
    InMux I__1614 (
            .O(N__7546),
            .I(N__7543));
    LocalMux I__1613 (
            .O(N__7543),
            .I(N__7540));
    Span4Mux_v I__1612 (
            .O(N__7540),
            .I(N__7537));
    Span4Mux_v I__1611 (
            .O(N__7537),
            .I(N__7534));
    Span4Mux_h I__1610 (
            .O(N__7534),
            .I(N__7530));
    IoInMux I__1609 (
            .O(N__7533),
            .I(N__7527));
    Odrv4 I__1608 (
            .O(N__7530),
            .I(CharacterDisplay__decfrac8));
    LocalMux I__1607 (
            .O(N__7527),
            .I(CharacterDisplay__decfrac8));
    InMux I__1606 (
            .O(N__7522),
            .I(N__7513));
    InMux I__1605 (
            .O(N__7521),
            .I(N__7513));
    InMux I__1604 (
            .O(N__7520),
            .I(N__7513));
    LocalMux I__1603 (
            .O(N__7513),
            .I(G_255));
    InMux I__1602 (
            .O(N__7510),
            .I(N__7501));
    InMux I__1601 (
            .O(N__7509),
            .I(N__7501));
    InMux I__1600 (
            .O(N__7508),
            .I(N__7501));
    LocalMux I__1599 (
            .O(N__7501),
            .I(G_254));
    CascadeMux I__1598 (
            .O(N__7498),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4_cascade_));
    InMux I__1597 (
            .O(N__7495),
            .I(N__7492));
    LocalMux I__1596 (
            .O(N__7492),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i_8));
    InMux I__1595 (
            .O(N__7489),
            .I(N__7485));
    InMux I__1594 (
            .O(N__7488),
            .I(N__7482));
    LocalMux I__1593 (
            .O(N__7485),
            .I(visibleXZ0Z_7));
    LocalMux I__1592 (
            .O(N__7482),
            .I(visibleXZ0Z_7));
    CascadeMux I__1591 (
            .O(N__7477),
            .I(N__7474));
    InMux I__1590 (
            .O(N__7474),
            .I(N__7471));
    LocalMux I__1589 (
            .O(N__7471),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i));
    InMux I__1588 (
            .O(N__7468),
            .I(N__7463));
    InMux I__1587 (
            .O(N__7467),
            .I(N__7460));
    CascadeMux I__1586 (
            .O(N__7466),
            .I(N__7451));
    LocalMux I__1585 (
            .O(N__7463),
            .I(N__7444));
    LocalMux I__1584 (
            .O(N__7460),
            .I(N__7444));
    InMux I__1583 (
            .O(N__7459),
            .I(N__7441));
    InMux I__1582 (
            .O(N__7458),
            .I(N__7423));
    InMux I__1581 (
            .O(N__7457),
            .I(N__7423));
    InMux I__1580 (
            .O(N__7456),
            .I(N__7423));
    InMux I__1579 (
            .O(N__7455),
            .I(N__7423));
    InMux I__1578 (
            .O(N__7454),
            .I(N__7423));
    InMux I__1577 (
            .O(N__7451),
            .I(N__7420));
    InMux I__1576 (
            .O(N__7450),
            .I(N__7415));
    InMux I__1575 (
            .O(N__7449),
            .I(N__7415));
    Span4Mux_v I__1574 (
            .O(N__7444),
            .I(N__7410));
    LocalMux I__1573 (
            .O(N__7441),
            .I(N__7410));
    InMux I__1572 (
            .O(N__7440),
            .I(N__7405));
    InMux I__1571 (
            .O(N__7439),
            .I(N__7405));
    InMux I__1570 (
            .O(N__7438),
            .I(N__7398));
    InMux I__1569 (
            .O(N__7437),
            .I(N__7398));
    InMux I__1568 (
            .O(N__7436),
            .I(N__7398));
    InMux I__1567 (
            .O(N__7435),
            .I(N__7395));
    InMux I__1566 (
            .O(N__7434),
            .I(N__7392));
    LocalMux I__1565 (
            .O(N__7423),
            .I(CO3_0));
    LocalMux I__1564 (
            .O(N__7420),
            .I(CO3_0));
    LocalMux I__1563 (
            .O(N__7415),
            .I(CO3_0));
    Odrv4 I__1562 (
            .O(N__7410),
            .I(CO3_0));
    LocalMux I__1561 (
            .O(N__7405),
            .I(CO3_0));
    LocalMux I__1560 (
            .O(N__7398),
            .I(CO3_0));
    LocalMux I__1559 (
            .O(N__7395),
            .I(CO3_0));
    LocalMux I__1558 (
            .O(N__7392),
            .I(CO3_0));
    ClkMux I__1557 (
            .O(N__7375),
            .I(N__7306));
    ClkMux I__1556 (
            .O(N__7374),
            .I(N__7306));
    ClkMux I__1555 (
            .O(N__7373),
            .I(N__7306));
    ClkMux I__1554 (
            .O(N__7372),
            .I(N__7306));
    ClkMux I__1553 (
            .O(N__7371),
            .I(N__7306));
    ClkMux I__1552 (
            .O(N__7370),
            .I(N__7306));
    ClkMux I__1551 (
            .O(N__7369),
            .I(N__7306));
    ClkMux I__1550 (
            .O(N__7368),
            .I(N__7306));
    ClkMux I__1549 (
            .O(N__7367),
            .I(N__7306));
    ClkMux I__1548 (
            .O(N__7366),
            .I(N__7306));
    ClkMux I__1547 (
            .O(N__7365),
            .I(N__7306));
    ClkMux I__1546 (
            .O(N__7364),
            .I(N__7306));
    ClkMux I__1545 (
            .O(N__7363),
            .I(N__7306));
    ClkMux I__1544 (
            .O(N__7362),
            .I(N__7306));
    ClkMux I__1543 (
            .O(N__7361),
            .I(N__7306));
    ClkMux I__1542 (
            .O(N__7360),
            .I(N__7306));
    ClkMux I__1541 (
            .O(N__7359),
            .I(N__7306));
    ClkMux I__1540 (
            .O(N__7358),
            .I(N__7306));
    ClkMux I__1539 (
            .O(N__7357),
            .I(N__7306));
    ClkMux I__1538 (
            .O(N__7356),
            .I(N__7306));
    ClkMux I__1537 (
            .O(N__7355),
            .I(N__7306));
    ClkMux I__1536 (
            .O(N__7354),
            .I(N__7306));
    ClkMux I__1535 (
            .O(N__7353),
            .I(N__7306));
    GlobalMux I__1534 (
            .O(N__7306),
            .I(N__7303));
    gio2CtrlBuf I__1533 (
            .O(N__7303),
            .I(PixelClock_g));
    CEMux I__1532 (
            .O(N__7300),
            .I(N__7258));
    CEMux I__1531 (
            .O(N__7299),
            .I(N__7258));
    CEMux I__1530 (
            .O(N__7298),
            .I(N__7258));
    CEMux I__1529 (
            .O(N__7297),
            .I(N__7258));
    CEMux I__1528 (
            .O(N__7296),
            .I(N__7258));
    CEMux I__1527 (
            .O(N__7295),
            .I(N__7258));
    CEMux I__1526 (
            .O(N__7294),
            .I(N__7258));
    CEMux I__1525 (
            .O(N__7293),
            .I(N__7258));
    CEMux I__1524 (
            .O(N__7292),
            .I(N__7258));
    CEMux I__1523 (
            .O(N__7291),
            .I(N__7258));
    CEMux I__1522 (
            .O(N__7290),
            .I(N__7258));
    CEMux I__1521 (
            .O(N__7289),
            .I(N__7258));
    CEMux I__1520 (
            .O(N__7288),
            .I(N__7258));
    CEMux I__1519 (
            .O(N__7287),
            .I(N__7258));
    GlobalMux I__1518 (
            .O(N__7258),
            .I(N__7255));
    gio2CtrlBuf I__1517 (
            .O(N__7255),
            .I(un15_beamy_g));
    CascadeMux I__1516 (
            .O(N__7252),
            .I(N__7249));
    InMux I__1515 (
            .O(N__7249),
            .I(N__7246));
    LocalMux I__1514 (
            .O(N__7246),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8PZ0Z8));
    InMux I__1513 (
            .O(N__7243),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    CascadeMux I__1512 (
            .O(N__7240),
            .I(N__7237));
    InMux I__1511 (
            .O(N__7237),
            .I(N__7234));
    LocalMux I__1510 (
            .O(N__7234),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQZ0Z8));
    InMux I__1509 (
            .O(N__7231),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__1508 (
            .O(N__7228),
            .I(N__7225));
    LocalMux I__1507 (
            .O(N__7225),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO));
    InMux I__1506 (
            .O(N__7222),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    InMux I__1505 (
            .O(N__7219),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7));
    InMux I__1504 (
            .O(N__7216),
            .I(N__7213));
    LocalMux I__1503 (
            .O(N__7213),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEAZ0Z08));
    InMux I__1502 (
            .O(N__7210),
            .I(N__7207));
    LocalMux I__1501 (
            .O(N__7207),
            .I(N__7201));
    CascadeMux I__1500 (
            .O(N__7206),
            .I(N__7198));
    InMux I__1499 (
            .O(N__7205),
            .I(N__7195));
    InMux I__1498 (
            .O(N__7204),
            .I(N__7192));
    Span4Mux_v I__1497 (
            .O(N__7201),
            .I(N__7189));
    InMux I__1496 (
            .O(N__7198),
            .I(N__7186));
    LocalMux I__1495 (
            .O(N__7195),
            .I(N__7183));
    LocalMux I__1494 (
            .O(N__7192),
            .I(beamXZ0Z_10));
    Odrv4 I__1493 (
            .O(N__7189),
            .I(beamXZ0Z_10));
    LocalMux I__1492 (
            .O(N__7186),
            .I(beamXZ0Z_10));
    Odrv4 I__1491 (
            .O(N__7183),
            .I(beamXZ0Z_10));
    InMux I__1490 (
            .O(N__7174),
            .I(N__7171));
    LocalMux I__1489 (
            .O(N__7171),
            .I(N__7168));
    Span4Mux_h I__1488 (
            .O(N__7168),
            .I(N__7162));
    InMux I__1487 (
            .O(N__7167),
            .I(N__7159));
    InMux I__1486 (
            .O(N__7166),
            .I(N__7154));
    InMux I__1485 (
            .O(N__7165),
            .I(N__7154));
    Odrv4 I__1484 (
            .O(N__7162),
            .I(un1_beamx_2));
    LocalMux I__1483 (
            .O(N__7159),
            .I(un1_beamx_2));
    LocalMux I__1482 (
            .O(N__7154),
            .I(un1_beamx_2));
    CascadeMux I__1481 (
            .O(N__7147),
            .I(N__7144));
    InMux I__1480 (
            .O(N__7144),
            .I(N__7141));
    LocalMux I__1479 (
            .O(N__7141),
            .I(N__7132));
    InMux I__1478 (
            .O(N__7140),
            .I(N__7129));
    InMux I__1477 (
            .O(N__7139),
            .I(N__7126));
    InMux I__1476 (
            .O(N__7138),
            .I(N__7119));
    InMux I__1475 (
            .O(N__7137),
            .I(N__7119));
    InMux I__1474 (
            .O(N__7136),
            .I(N__7119));
    InMux I__1473 (
            .O(N__7135),
            .I(N__7116));
    Odrv12 I__1472 (
            .O(N__7132),
            .I(beamXZ0Z_7));
    LocalMux I__1471 (
            .O(N__7129),
            .I(beamXZ0Z_7));
    LocalMux I__1470 (
            .O(N__7126),
            .I(beamXZ0Z_7));
    LocalMux I__1469 (
            .O(N__7119),
            .I(beamXZ0Z_7));
    LocalMux I__1468 (
            .O(N__7116),
            .I(beamXZ0Z_7));
    InMux I__1467 (
            .O(N__7105),
            .I(N__7102));
    LocalMux I__1466 (
            .O(N__7102),
            .I(un1_beamxlt10_0));
    IoInMux I__1465 (
            .O(N__7099),
            .I(N__7096));
    LocalMux I__1464 (
            .O(N__7096),
            .I(N__7093));
    IoSpan4Mux I__1463 (
            .O(N__7093),
            .I(N__7089));
    IoInMux I__1462 (
            .O(N__7092),
            .I(N__7086));
    Span4Mux_s2_v I__1461 (
            .O(N__7089),
            .I(N__7083));
    LocalMux I__1460 (
            .O(N__7086),
            .I(N__7080));
    Sp12to4 I__1459 (
            .O(N__7083),
            .I(N__7075));
    Span12Mux_s1_v I__1458 (
            .O(N__7080),
            .I(N__7075));
    Odrv12 I__1457 (
            .O(N__7075),
            .I(HSync_c));
    CascadeMux I__1456 (
            .O(N__7072),
            .I(N__7069));
    InMux I__1455 (
            .O(N__7069),
            .I(N__7066));
    LocalMux I__1454 (
            .O(N__7066),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i));
    InMux I__1453 (
            .O(N__7063),
            .I(N__7059));
    InMux I__1452 (
            .O(N__7062),
            .I(N__7056));
    LocalMux I__1451 (
            .O(N__7059),
            .I(visibleXZ0Z_6));
    LocalMux I__1450 (
            .O(N__7056),
            .I(visibleXZ0Z_6));
    InMux I__1449 (
            .O(N__7051),
            .I(N__7048));
    LocalMux I__1448 (
            .O(N__7048),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTKZ0Z2));
    InMux I__1447 (
            .O(N__7045),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__1446 (
            .O(N__7042),
            .I(N__7038));
    InMux I__1445 (
            .O(N__7041),
            .I(N__7035));
    LocalMux I__1444 (
            .O(N__7038),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412));
    LocalMux I__1443 (
            .O(N__7035),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412));
    CascadeMux I__1442 (
            .O(N__7030),
            .I(N__7027));
    InMux I__1441 (
            .O(N__7027),
            .I(N__7024));
    LocalMux I__1440 (
            .O(N__7024),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BDZ0Z1));
    CascadeMux I__1439 (
            .O(N__7021),
            .I(N__7017));
    InMux I__1438 (
            .O(N__7020),
            .I(N__7012));
    InMux I__1437 (
            .O(N__7017),
            .I(N__7012));
    LocalMux I__1436 (
            .O(N__7012),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19MZ0Z3));
    InMux I__1435 (
            .O(N__7009),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__1434 (
            .O(N__7006),
            .I(N__7000));
    InMux I__1433 (
            .O(N__7005),
            .I(N__7000));
    LocalMux I__1432 (
            .O(N__7000),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i_8));
    CascadeMux I__1431 (
            .O(N__6997),
            .I(N__6994));
    InMux I__1430 (
            .O(N__6994),
            .I(N__6991));
    LocalMux I__1429 (
            .O(N__6991),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMKZ0Z642));
    InMux I__1428 (
            .O(N__6988),
            .I(N__6985));
    LocalMux I__1427 (
            .O(N__6985),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_axb_8));
    InMux I__1426 (
            .O(N__6982),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    InMux I__1425 (
            .O(N__6979),
            .I(N__6976));
    LocalMux I__1424 (
            .O(N__6976),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_axb_8));
    InMux I__1423 (
            .O(N__6973),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7));
    CascadeMux I__1422 (
            .O(N__6970),
            .I(N__6966));
    InMux I__1421 (
            .O(N__6969),
            .I(N__6962));
    InMux I__1420 (
            .O(N__6966),
            .I(N__6957));
    InMux I__1419 (
            .O(N__6965),
            .I(N__6957));
    LocalMux I__1418 (
            .O(N__6962),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4));
    LocalMux I__1417 (
            .O(N__6957),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4));
    CascadeMux I__1416 (
            .O(N__6952),
            .I(N__6949));
    InMux I__1415 (
            .O(N__6949),
            .I(N__6946));
    LocalMux I__1414 (
            .O(N__6946),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKVZ0));
    InMux I__1413 (
            .O(N__6943),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__1412 (
            .O(N__6940),
            .I(N__6937));
    LocalMux I__1411 (
            .O(N__6937),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_axb_8));
    InMux I__1410 (
            .O(N__6934),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__1409 (
            .O(N__6931),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7));
    InMux I__1408 (
            .O(N__6928),
            .I(N__6923));
    InMux I__1407 (
            .O(N__6927),
            .I(N__6918));
    InMux I__1406 (
            .O(N__6926),
            .I(N__6918));
    LocalMux I__1405 (
            .O(N__6923),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0));
    LocalMux I__1404 (
            .O(N__6918),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0));
    InMux I__1403 (
            .O(N__6913),
            .I(N__6907));
    InMux I__1402 (
            .O(N__6912),
            .I(N__6907));
    LocalMux I__1401 (
            .O(N__6907),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i_8));
    InMux I__1400 (
            .O(N__6904),
            .I(N__6900));
    InMux I__1399 (
            .O(N__6903),
            .I(N__6897));
    LocalMux I__1398 (
            .O(N__6900),
            .I(N__6892));
    LocalMux I__1397 (
            .O(N__6897),
            .I(N__6892));
    Span4Mux_h I__1396 (
            .O(N__6892),
            .I(N__6889));
    Odrv4 I__1395 (
            .O(N__6889),
            .I(visibleXZ0Z_5));
    InMux I__1394 (
            .O(N__6886),
            .I(N__6883));
    LocalMux I__1393 (
            .O(N__6883),
            .I(N__6880));
    Odrv4 I__1392 (
            .O(N__6880),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56BZ0Z05));
    InMux I__1391 (
            .O(N__6877),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__1390 (
            .O(N__6874),
            .I(N__6871));
    InMux I__1389 (
            .O(N__6871),
            .I(N__6868));
    LocalMux I__1388 (
            .O(N__6868),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNICZ0Z7997));
    InMux I__1387 (
            .O(N__6865),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__1386 (
            .O(N__6862),
            .I(N__6859));
    LocalMux I__1385 (
            .O(N__6859),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_axb_8));
    InMux I__1384 (
            .O(N__6856),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__1383 (
            .O(N__6853),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7));
    CascadeMux I__1382 (
            .O(N__6850),
            .I(N__6846));
    InMux I__1381 (
            .O(N__6849),
            .I(N__6842));
    InMux I__1380 (
            .O(N__6846),
            .I(N__6837));
    InMux I__1379 (
            .O(N__6845),
            .I(N__6837));
    LocalMux I__1378 (
            .O(N__6842),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19));
    LocalMux I__1377 (
            .O(N__6837),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19));
    InMux I__1376 (
            .O(N__6832),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__1375 (
            .O(N__6829),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__1374 (
            .O(N__6826),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    InMux I__1373 (
            .O(N__6823),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7));
    CascadeMux I__1372 (
            .O(N__6820),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412_cascade_));
    CascadeMux I__1371 (
            .O(N__6817),
            .I(N__6814));
    InMux I__1370 (
            .O(N__6814),
            .I(N__6811));
    LocalMux I__1369 (
            .O(N__6811),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i));
    InMux I__1368 (
            .O(N__6808),
            .I(N__6804));
    InMux I__1367 (
            .O(N__6807),
            .I(N__6797));
    LocalMux I__1366 (
            .O(N__6804),
            .I(N__6794));
    InMux I__1365 (
            .O(N__6803),
            .I(N__6785));
    InMux I__1364 (
            .O(N__6802),
            .I(N__6785));
    InMux I__1363 (
            .O(N__6801),
            .I(N__6785));
    InMux I__1362 (
            .O(N__6800),
            .I(N__6785));
    LocalMux I__1361 (
            .O(N__6797),
            .I(N_3_0));
    Odrv4 I__1360 (
            .O(N__6794),
            .I(N_3_0));
    LocalMux I__1359 (
            .O(N__6785),
            .I(N_3_0));
    InMux I__1358 (
            .O(N__6778),
            .I(N__6775));
    LocalMux I__1357 (
            .O(N__6775),
            .I(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx));
    InMux I__1356 (
            .O(N__6772),
            .I(N__6768));
    InMux I__1355 (
            .O(N__6771),
            .I(N__6765));
    LocalMux I__1354 (
            .O(N__6768),
            .I(visibleXZ0Z_8));
    LocalMux I__1353 (
            .O(N__6765),
            .I(visibleXZ0Z_8));
    CascadeMux I__1352 (
            .O(N__6760),
            .I(N__6757));
    InMux I__1351 (
            .O(N__6757),
            .I(N__6754));
    LocalMux I__1350 (
            .O(N__6754),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29RZ0Z21));
    InMux I__1349 (
            .O(N__6751),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    CascadeMux I__1348 (
            .O(N__6748),
            .I(N__6740));
    InMux I__1347 (
            .O(N__6747),
            .I(N__6737));
    InMux I__1346 (
            .O(N__6746),
            .I(N__6732));
    InMux I__1345 (
            .O(N__6745),
            .I(N__6732));
    InMux I__1344 (
            .O(N__6744),
            .I(N__6727));
    InMux I__1343 (
            .O(N__6743),
            .I(N__6727));
    InMux I__1342 (
            .O(N__6740),
            .I(N__6724));
    LocalMux I__1341 (
            .O(N__6737),
            .I(beamXZ0Z_6));
    LocalMux I__1340 (
            .O(N__6732),
            .I(beamXZ0Z_6));
    LocalMux I__1339 (
            .O(N__6727),
            .I(beamXZ0Z_6));
    LocalMux I__1338 (
            .O(N__6724),
            .I(beamXZ0Z_6));
    InMux I__1337 (
            .O(N__6715),
            .I(N__6707));
    InMux I__1336 (
            .O(N__6714),
            .I(N__6702));
    InMux I__1335 (
            .O(N__6713),
            .I(N__6702));
    InMux I__1334 (
            .O(N__6712),
            .I(N__6697));
    InMux I__1333 (
            .O(N__6711),
            .I(N__6697));
    InMux I__1332 (
            .O(N__6710),
            .I(N__6694));
    LocalMux I__1331 (
            .O(N__6707),
            .I(beamXZ0Z_4));
    LocalMux I__1330 (
            .O(N__6702),
            .I(beamXZ0Z_4));
    LocalMux I__1329 (
            .O(N__6697),
            .I(beamXZ0Z_4));
    LocalMux I__1328 (
            .O(N__6694),
            .I(beamXZ0Z_4));
    CascadeMux I__1327 (
            .O(N__6685),
            .I(N__6680));
    CascadeMux I__1326 (
            .O(N__6684),
            .I(N__6675));
    InMux I__1325 (
            .O(N__6683),
            .I(N__6671));
    InMux I__1324 (
            .O(N__6680),
            .I(N__6666));
    InMux I__1323 (
            .O(N__6679),
            .I(N__6666));
    InMux I__1322 (
            .O(N__6678),
            .I(N__6661));
    InMux I__1321 (
            .O(N__6675),
            .I(N__6661));
    InMux I__1320 (
            .O(N__6674),
            .I(N__6658));
    LocalMux I__1319 (
            .O(N__6671),
            .I(beamXZ0Z_5));
    LocalMux I__1318 (
            .O(N__6666),
            .I(beamXZ0Z_5));
    LocalMux I__1317 (
            .O(N__6661),
            .I(beamXZ0Z_5));
    LocalMux I__1316 (
            .O(N__6658),
            .I(beamXZ0Z_5));
    CascadeMux I__1315 (
            .O(N__6649),
            .I(N__6643));
    InMux I__1314 (
            .O(N__6648),
            .I(N__6639));
    InMux I__1313 (
            .O(N__6647),
            .I(N__6634));
    InMux I__1312 (
            .O(N__6646),
            .I(N__6634));
    InMux I__1311 (
            .O(N__6643),
            .I(N__6631));
    InMux I__1310 (
            .O(N__6642),
            .I(N__6628));
    LocalMux I__1309 (
            .O(N__6639),
            .I(beamXZ0Z_3));
    LocalMux I__1308 (
            .O(N__6634),
            .I(beamXZ0Z_3));
    LocalMux I__1307 (
            .O(N__6631),
            .I(beamXZ0Z_3));
    LocalMux I__1306 (
            .O(N__6628),
            .I(beamXZ0Z_3));
    InMux I__1305 (
            .O(N__6619),
            .I(N__6611));
    InMux I__1304 (
            .O(N__6618),
            .I(N__6611));
    InMux I__1303 (
            .O(N__6617),
            .I(N__6605));
    InMux I__1302 (
            .O(N__6616),
            .I(N__6605));
    LocalMux I__1301 (
            .O(N__6611),
            .I(N__6602));
    InMux I__1300 (
            .O(N__6610),
            .I(N__6599));
    LocalMux I__1299 (
            .O(N__6605),
            .I(N__6596));
    Odrv4 I__1298 (
            .O(N__6602),
            .I(c_if_generate_plus_mult1_un47_sum_1));
    LocalMux I__1297 (
            .O(N__6599),
            .I(c_if_generate_plus_mult1_un47_sum_1));
    Odrv4 I__1296 (
            .O(N__6596),
            .I(c_if_generate_plus_mult1_un47_sum_1));
    InMux I__1295 (
            .O(N__6589),
            .I(N__6586));
    LocalMux I__1294 (
            .O(N__6586),
            .I(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx));
    CascadeMux I__1293 (
            .O(N__6583),
            .I(N__6580));
    InMux I__1292 (
            .O(N__6580),
            .I(N__6577));
    LocalMux I__1291 (
            .O(N__6577),
            .I(un5_vx_i_25));
    InMux I__1290 (
            .O(N__6574),
            .I(N__6571));
    LocalMux I__1289 (
            .O(N__6571),
            .I(N__6568));
    Span4Mux_h I__1288 (
            .O(N__6568),
            .I(N__6565));
    Odrv4 I__1287 (
            .O(N__6565),
            .I(c_if_generate_plus_mult1_un47_sum0_2));
    InMux I__1286 (
            .O(N__6562),
            .I(c_if_generate_plus_mult1_un47_sum_0_cry_1));
    InMux I__1285 (
            .O(N__6559),
            .I(N__6556));
    LocalMux I__1284 (
            .O(N__6556),
            .I(if_generate_plus_mult1_un47_sum_0_cry_3_ma));
    CascadeMux I__1283 (
            .O(N__6553),
            .I(N__6550));
    InMux I__1282 (
            .O(N__6550),
            .I(N__6547));
    LocalMux I__1281 (
            .O(N__6547),
            .I(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx));
    InMux I__1280 (
            .O(N__6544),
            .I(N__6541));
    LocalMux I__1279 (
            .O(N__6541),
            .I(N__6538));
    Odrv4 I__1278 (
            .O(N__6538),
            .I(c_if_generate_plus_mult1_un47_sum0_3));
    InMux I__1277 (
            .O(N__6535),
            .I(c_if_generate_plus_mult1_un47_sum_0_cry_2));
    CascadeMux I__1276 (
            .O(N__6532),
            .I(N__6529));
    InMux I__1275 (
            .O(N__6529),
            .I(N__6526));
    LocalMux I__1274 (
            .O(N__6526),
            .I(N_186_0_i));
    InMux I__1273 (
            .O(N__6523),
            .I(N__6520));
    LocalMux I__1272 (
            .O(N__6520),
            .I(N__6517));
    Odrv4 I__1271 (
            .O(N__6517),
            .I(c_if_generate_plus_mult1_un47_sum0_4));
    InMux I__1270 (
            .O(N__6514),
            .I(c_if_generate_plus_mult1_un47_sum_0_cry_3));
    InMux I__1269 (
            .O(N__6511),
            .I(c_if_generate_plus_mult1_un47_sum_0_cry_4));
    InMux I__1268 (
            .O(N__6508),
            .I(N__6505));
    LocalMux I__1267 (
            .O(N__6505),
            .I(N__6500));
    InMux I__1266 (
            .O(N__6504),
            .I(N__6495));
    InMux I__1265 (
            .O(N__6503),
            .I(N__6495));
    Span4Mux_v I__1264 (
            .O(N__6500),
            .I(N__6492));
    LocalMux I__1263 (
            .O(N__6495),
            .I(N__6489));
    Odrv4 I__1262 (
            .O(N__6492),
            .I(c_if_generate_plus_mult1_un47_sum0_5));
    Odrv4 I__1261 (
            .O(N__6489),
            .I(c_if_generate_plus_mult1_un47_sum0_5));
    InMux I__1260 (
            .O(N__6484),
            .I(N__6481));
    LocalMux I__1259 (
            .O(N__6481),
            .I(N__6471));
    InMux I__1258 (
            .O(N__6480),
            .I(N__6468));
    InMux I__1257 (
            .O(N__6479),
            .I(N__6465));
    InMux I__1256 (
            .O(N__6478),
            .I(N__6460));
    InMux I__1255 (
            .O(N__6477),
            .I(N__6460));
    InMux I__1254 (
            .O(N__6476),
            .I(N__6453));
    InMux I__1253 (
            .O(N__6475),
            .I(N__6453));
    InMux I__1252 (
            .O(N__6474),
            .I(N__6453));
    Odrv4 I__1251 (
            .O(N__6471),
            .I(un5_vx_cry_6_c_RNI59BZ0));
    LocalMux I__1250 (
            .O(N__6468),
            .I(un5_vx_cry_6_c_RNI59BZ0));
    LocalMux I__1249 (
            .O(N__6465),
            .I(un5_vx_cry_6_c_RNI59BZ0));
    LocalMux I__1248 (
            .O(N__6460),
            .I(un5_vx_cry_6_c_RNI59BZ0));
    LocalMux I__1247 (
            .O(N__6453),
            .I(un5_vx_cry_6_c_RNI59BZ0));
    InMux I__1246 (
            .O(N__6442),
            .I(N__6436));
    InMux I__1245 (
            .O(N__6441),
            .I(N__6436));
    LocalMux I__1244 (
            .O(N__6436),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i_8));
    InMux I__1243 (
            .O(N__6433),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7));
    InMux I__1242 (
            .O(N__6430),
            .I(N__6427));
    LocalMux I__1241 (
            .O(N__6427),
            .I(N__6424));
    Span4Mux_h I__1240 (
            .O(N__6424),
            .I(N__6421));
    Odrv4 I__1239 (
            .O(N__6421),
            .I(N_84));
    CascadeMux I__1238 (
            .O(N__6418),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0_cascade_));
    InMux I__1237 (
            .O(N__6415),
            .I(N__6412));
    LocalMux I__1236 (
            .O(N__6412),
            .I(N_53));
    InMux I__1235 (
            .O(N__6409),
            .I(N__6405));
    InMux I__1234 (
            .O(N__6408),
            .I(N__6402));
    LocalMux I__1233 (
            .O(N__6405),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0));
    LocalMux I__1232 (
            .O(N__6402),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0));
    InMux I__1231 (
            .O(N__6397),
            .I(N__6394));
    LocalMux I__1230 (
            .O(N__6394),
            .I(Pixel_RNOZ0Z_8));
    CascadeMux I__1229 (
            .O(N__6391),
            .I(N__6388));
    InMux I__1228 (
            .O(N__6388),
            .I(N__6379));
    InMux I__1227 (
            .O(N__6387),
            .I(N__6379));
    InMux I__1226 (
            .O(N__6386),
            .I(N__6379));
    LocalMux I__1225 (
            .O(N__6379),
            .I(N__6376));
    Span4Mux_v I__1224 (
            .O(N__6376),
            .I(N__6373));
    Span4Mux_h I__1223 (
            .O(N__6373),
            .I(N__6370));
    Odrv4 I__1222 (
            .O(N__6370),
            .I(visibleXZ0Z_4));
    InMux I__1221 (
            .O(N__6367),
            .I(N__6364));
    LocalMux I__1220 (
            .O(N__6364),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0));
    InMux I__1219 (
            .O(N__6361),
            .I(N__6358));
    LocalMux I__1218 (
            .O(N__6358),
            .I(N_81));
    CascadeMux I__1217 (
            .O(N__6355),
            .I(N__6352));
    InMux I__1216 (
            .O(N__6352),
            .I(N__6349));
    LocalMux I__1215 (
            .O(N__6349),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i));
    InMux I__1214 (
            .O(N__6346),
            .I(N__6340));
    InMux I__1213 (
            .O(N__6345),
            .I(N__6337));
    InMux I__1212 (
            .O(N__6344),
            .I(N__6334));
    InMux I__1211 (
            .O(N__6343),
            .I(N__6331));
    LocalMux I__1210 (
            .O(N__6340),
            .I(beamXZ0Z_2));
    LocalMux I__1209 (
            .O(N__6337),
            .I(beamXZ0Z_2));
    LocalMux I__1208 (
            .O(N__6334),
            .I(beamXZ0Z_2));
    LocalMux I__1207 (
            .O(N__6331),
            .I(beamXZ0Z_2));
    InMux I__1206 (
            .O(N__6322),
            .I(N__6319));
    LocalMux I__1205 (
            .O(N__6319),
            .I(N__6315));
    InMux I__1204 (
            .O(N__6318),
            .I(N__6310));
    Span4Mux_v I__1203 (
            .O(N__6315),
            .I(N__6307));
    InMux I__1202 (
            .O(N__6314),
            .I(N__6304));
    InMux I__1201 (
            .O(N__6313),
            .I(N__6301));
    LocalMux I__1200 (
            .O(N__6310),
            .I(beamXZ0Z_1));
    Odrv4 I__1199 (
            .O(N__6307),
            .I(beamXZ0Z_1));
    LocalMux I__1198 (
            .O(N__6304),
            .I(beamXZ0Z_1));
    LocalMux I__1197 (
            .O(N__6301),
            .I(beamXZ0Z_1));
    CascadeMux I__1196 (
            .O(N__6292),
            .I(un3_beamx_5_cascade_));
    CascadeMux I__1195 (
            .O(N__6289),
            .I(N__6285));
    InMux I__1194 (
            .O(N__6288),
            .I(N__6278));
    InMux I__1193 (
            .O(N__6285),
            .I(N__6275));
    InMux I__1192 (
            .O(N__6284),
            .I(N__6272));
    InMux I__1191 (
            .O(N__6283),
            .I(N__6269));
    InMux I__1190 (
            .O(N__6282),
            .I(N__6264));
    InMux I__1189 (
            .O(N__6281),
            .I(N__6264));
    LocalMux I__1188 (
            .O(N__6278),
            .I(un5_vx));
    LocalMux I__1187 (
            .O(N__6275),
            .I(un5_vx));
    LocalMux I__1186 (
            .O(N__6272),
            .I(un5_vx));
    LocalMux I__1185 (
            .O(N__6269),
            .I(un5_vx));
    LocalMux I__1184 (
            .O(N__6264),
            .I(un5_vx));
    CascadeMux I__1183 (
            .O(N__6253),
            .I(un3_beamx_7_cascade_));
    CEMux I__1182 (
            .O(N__6250),
            .I(N__6245));
    InMux I__1181 (
            .O(N__6249),
            .I(N__6240));
    InMux I__1180 (
            .O(N__6248),
            .I(N__6240));
    LocalMux I__1179 (
            .O(N__6245),
            .I(N__6236));
    LocalMux I__1178 (
            .O(N__6240),
            .I(N__6231));
    InMux I__1177 (
            .O(N__6239),
            .I(N__6228));
    Span4Mux_h I__1176 (
            .O(N__6236),
            .I(N__6225));
    InMux I__1175 (
            .O(N__6235),
            .I(N__6220));
    InMux I__1174 (
            .O(N__6234),
            .I(N__6220));
    Span4Mux_v I__1173 (
            .O(N__6231),
            .I(N__6217));
    LocalMux I__1172 (
            .O(N__6228),
            .I(N__6212));
    Span4Mux_v I__1171 (
            .O(N__6225),
            .I(N__6212));
    LocalMux I__1170 (
            .O(N__6220),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__1169 (
            .O(N__6217),
            .I(beamX_RNI5457Z0Z_5));
    Odrv4 I__1168 (
            .O(N__6212),
            .I(beamX_RNI5457Z0Z_5));
    CascadeMux I__1167 (
            .O(N__6205),
            .I(N__6202));
    InMux I__1166 (
            .O(N__6202),
            .I(N__6199));
    LocalMux I__1165 (
            .O(N__6199),
            .I(if_generate_plus_mult1_un54_sum_axb_2_l_fx));
    CascadeMux I__1164 (
            .O(N__6196),
            .I(N__6193));
    InMux I__1163 (
            .O(N__6193),
            .I(N__6190));
    LocalMux I__1162 (
            .O(N__6190),
            .I(N__6187));
    Odrv4 I__1161 (
            .O(N__6187),
            .I(if_generate_plus_mult1_un54_sum_cry_2_s));
    InMux I__1160 (
            .O(N__6184),
            .I(c_if_generate_plus_mult1_un54_sum_cry_1));
    InMux I__1159 (
            .O(N__6181),
            .I(N__6178));
    LocalMux I__1158 (
            .O(N__6178),
            .I(if_generate_plus_mult1_un54_sum_axb_3_l_fx));
    CascadeMux I__1157 (
            .O(N__6175),
            .I(N__6172));
    InMux I__1156 (
            .O(N__6172),
            .I(N__6168));
    InMux I__1155 (
            .O(N__6171),
            .I(N__6165));
    LocalMux I__1154 (
            .O(N__6168),
            .I(N__6162));
    LocalMux I__1153 (
            .O(N__6165),
            .I(if_generate_plus_mult1_un47_sum_m_2));
    Odrv4 I__1152 (
            .O(N__6162),
            .I(if_generate_plus_mult1_un47_sum_m_2));
    CascadeMux I__1151 (
            .O(N__6157),
            .I(N__6154));
    InMux I__1150 (
            .O(N__6154),
            .I(N__6151));
    LocalMux I__1149 (
            .O(N__6151),
            .I(N__6148));
    Odrv4 I__1148 (
            .O(N__6148),
            .I(if_generate_plus_mult1_un54_sum_cry_3_s));
    InMux I__1147 (
            .O(N__6145),
            .I(c_if_generate_plus_mult1_un54_sum_cry_2));
    CascadeMux I__1146 (
            .O(N__6142),
            .I(N__6138));
    CascadeMux I__1145 (
            .O(N__6141),
            .I(N__6135));
    InMux I__1144 (
            .O(N__6138),
            .I(N__6130));
    InMux I__1143 (
            .O(N__6135),
            .I(N__6127));
    InMux I__1142 (
            .O(N__6134),
            .I(N__6122));
    InMux I__1141 (
            .O(N__6133),
            .I(N__6122));
    LocalMux I__1140 (
            .O(N__6130),
            .I(N_18));
    LocalMux I__1139 (
            .O(N__6127),
            .I(N_18));
    LocalMux I__1138 (
            .O(N__6122),
            .I(N_18));
    CascadeMux I__1137 (
            .O(N__6115),
            .I(N__6112));
    InMux I__1136 (
            .O(N__6112),
            .I(N__6109));
    LocalMux I__1135 (
            .O(N__6109),
            .I(if_generate_plus_mult1_un54_sum_axb_4_l_fx));
    InMux I__1134 (
            .O(N__6106),
            .I(N__6103));
    LocalMux I__1133 (
            .O(N__6103),
            .I(N__6100));
    Odrv4 I__1132 (
            .O(N__6100),
            .I(c_if_generate_plus_mult1_un61_sum_axbZ0Z_5));
    InMux I__1131 (
            .O(N__6097),
            .I(c_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__1130 (
            .O(N__6094),
            .I(N__6091));
    LocalMux I__1129 (
            .O(N__6091),
            .I(c_if_generate_plus_mult1_un54_sum_axbZ0Z_5));
    InMux I__1128 (
            .O(N__6088),
            .I(c_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__1127 (
            .O(N__6085),
            .I(N__6082));
    LocalMux I__1126 (
            .O(N__6082),
            .I(N__6079));
    Span4Mux_v I__1125 (
            .O(N__6079),
            .I(N__6075));
    InMux I__1124 (
            .O(N__6078),
            .I(N__6072));
    Span4Mux_v I__1123 (
            .O(N__6075),
            .I(N__6065));
    LocalMux I__1122 (
            .O(N__6072),
            .I(N__6065));
    InMux I__1121 (
            .O(N__6071),
            .I(N__6062));
    InMux I__1120 (
            .O(N__6070),
            .I(N__6059));
    Odrv4 I__1119 (
            .O(N__6065),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__1118 (
            .O(N__6062),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    LocalMux I__1117 (
            .O(N__6059),
            .I(if_generate_plus_mult1_un54_sum_s_5));
    InMux I__1116 (
            .O(N__6052),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__1115 (
            .O(N__6049),
            .I(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5));
    InMux I__1114 (
            .O(N__6046),
            .I(N__6043));
    LocalMux I__1113 (
            .O(N__6043),
            .I(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx));
    InMux I__1112 (
            .O(N__6040),
            .I(c_if_generate_plus_mult1_un47_sum_1_cry_3));
    InMux I__1111 (
            .O(N__6037),
            .I(c_if_generate_plus_mult1_un47_sum_1_cry_4));
    CascadeMux I__1110 (
            .O(N__6034),
            .I(N__6030));
    InMux I__1109 (
            .O(N__6033),
            .I(N__6021));
    InMux I__1108 (
            .O(N__6030),
            .I(N__6021));
    InMux I__1107 (
            .O(N__6029),
            .I(N__6018));
    InMux I__1106 (
            .O(N__6028),
            .I(N__6011));
    InMux I__1105 (
            .O(N__6027),
            .I(N__6011));
    InMux I__1104 (
            .O(N__6026),
            .I(N__6011));
    LocalMux I__1103 (
            .O(N__6021),
            .I(c_if_generate_plus_mult1_un47_sum_0_0));
    LocalMux I__1102 (
            .O(N__6018),
            .I(c_if_generate_plus_mult1_un47_sum_0_0));
    LocalMux I__1101 (
            .O(N__6011),
            .I(c_if_generate_plus_mult1_un47_sum_0_0));
    InMux I__1100 (
            .O(N__6004),
            .I(N__6001));
    LocalMux I__1099 (
            .O(N__6001),
            .I(c_if_generate_plus_mult1_un47_sum1_4));
    CascadeMux I__1098 (
            .O(N__5998),
            .I(N_18_cascade_));
    InMux I__1097 (
            .O(N__5995),
            .I(N__5992));
    LocalMux I__1096 (
            .O(N__5992),
            .I(c_if_generate_plus_mult1_un47_sum1_3));
    CascadeMux I__1095 (
            .O(N__5989),
            .I(N__5985));
    InMux I__1094 (
            .O(N__5988),
            .I(N__5981));
    InMux I__1093 (
            .O(N__5985),
            .I(N__5976));
    InMux I__1092 (
            .O(N__5984),
            .I(N__5976));
    LocalMux I__1091 (
            .O(N__5981),
            .I(c_if_generate_plus_mult1_un47_sum1_5));
    LocalMux I__1090 (
            .O(N__5976),
            .I(c_if_generate_plus_mult1_un47_sum1_5));
    InMux I__1089 (
            .O(N__5971),
            .I(N__5966));
    InMux I__1088 (
            .O(N__5970),
            .I(N__5961));
    InMux I__1087 (
            .O(N__5969),
            .I(N__5961));
    LocalMux I__1086 (
            .O(N__5966),
            .I(N__5956));
    LocalMux I__1085 (
            .O(N__5961),
            .I(N__5956));
    Odrv4 I__1084 (
            .O(N__5956),
            .I(c_if_generate_plus_mult1_un47_sum1_0));
    InMux I__1083 (
            .O(N__5953),
            .I(un8_beamx_cry_9));
    CascadeMux I__1082 (
            .O(N__5950),
            .I(un5_vx_i_25_cascade_));
    CascadeMux I__1081 (
            .O(N__5947),
            .I(N__5944));
    InMux I__1080 (
            .O(N__5944),
            .I(N__5941));
    LocalMux I__1079 (
            .O(N__5941),
            .I(un5_vx_i_0_25));
    InMux I__1078 (
            .O(N__5938),
            .I(c_if_generate_plus_mult1_un47_sum_1_cry_1));
    InMux I__1077 (
            .O(N__5935),
            .I(N__5932));
    LocalMux I__1076 (
            .O(N__5932),
            .I(c_if_generate_plus_mult1_un47_sum_0_axb_5_i));
    CascadeMux I__1075 (
            .O(N__5929),
            .I(N__5926));
    InMux I__1074 (
            .O(N__5926),
            .I(N__5923));
    LocalMux I__1073 (
            .O(N__5923),
            .I(N_13_0_i));
    InMux I__1072 (
            .O(N__5920),
            .I(c_if_generate_plus_mult1_un47_sum_1_cry_2));
    InMux I__1071 (
            .O(N__5917),
            .I(un8_beamx_cry_1));
    InMux I__1070 (
            .O(N__5914),
            .I(un8_beamx_cry_2));
    InMux I__1069 (
            .O(N__5911),
            .I(un8_beamx_cry_3));
    InMux I__1068 (
            .O(N__5908),
            .I(un8_beamx_cry_4));
    InMux I__1067 (
            .O(N__5905),
            .I(un8_beamx_cry_5));
    InMux I__1066 (
            .O(N__5902),
            .I(un8_beamx_cry_6));
    InMux I__1065 (
            .O(N__5899),
            .I(N__5893));
    InMux I__1064 (
            .O(N__5898),
            .I(N__5890));
    InMux I__1063 (
            .O(N__5897),
            .I(N__5885));
    InMux I__1062 (
            .O(N__5896),
            .I(N__5885));
    LocalMux I__1061 (
            .O(N__5893),
            .I(N__5882));
    LocalMux I__1060 (
            .O(N__5890),
            .I(beamXZ0Z_8));
    LocalMux I__1059 (
            .O(N__5885),
            .I(beamXZ0Z_8));
    Odrv4 I__1058 (
            .O(N__5882),
            .I(beamXZ0Z_8));
    InMux I__1057 (
            .O(N__5875),
            .I(un8_beamx_cry_7));
    CascadeMux I__1056 (
            .O(N__5872),
            .I(N__5868));
    InMux I__1055 (
            .O(N__5871),
            .I(N__5862));
    InMux I__1054 (
            .O(N__5868),
            .I(N__5862));
    InMux I__1053 (
            .O(N__5867),
            .I(N__5858));
    LocalMux I__1052 (
            .O(N__5862),
            .I(N__5855));
    InMux I__1051 (
            .O(N__5861),
            .I(N__5852));
    LocalMux I__1050 (
            .O(N__5858),
            .I(beamXZ0Z_9));
    Odrv4 I__1049 (
            .O(N__5855),
            .I(beamXZ0Z_9));
    LocalMux I__1048 (
            .O(N__5852),
            .I(beamXZ0Z_9));
    InMux I__1047 (
            .O(N__5845),
            .I(bfn_7_9_0_));
    InMux I__1046 (
            .O(N__5842),
            .I(N__5837));
    InMux I__1045 (
            .O(N__5841),
            .I(N__5832));
    InMux I__1044 (
            .O(N__5840),
            .I(N__5832));
    LocalMux I__1043 (
            .O(N__5837),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0));
    LocalMux I__1042 (
            .O(N__5832),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0));
    CascadeMux I__1041 (
            .O(N__5827),
            .I(N__5824));
    InMux I__1040 (
            .O(N__5824),
            .I(N__5818));
    InMux I__1039 (
            .O(N__5823),
            .I(N__5818));
    LocalMux I__1038 (
            .O(N__5818),
            .I(N__5815));
    Span4Mux_v I__1037 (
            .O(N__5815),
            .I(N__5812));
    Odrv4 I__1036 (
            .O(N__5812),
            .I(visibleYZ0Z_1));
    CascadeMux I__1035 (
            .O(N__5809),
            .I(N__5803));
    InMux I__1034 (
            .O(N__5808),
            .I(N__5798));
    InMux I__1033 (
            .O(N__5807),
            .I(N__5798));
    InMux I__1032 (
            .O(N__5806),
            .I(N__5795));
    InMux I__1031 (
            .O(N__5803),
            .I(N__5792));
    LocalMux I__1030 (
            .O(N__5798),
            .I(N__5789));
    LocalMux I__1029 (
            .O(N__5795),
            .I(visibleYZ0Z_2));
    LocalMux I__1028 (
            .O(N__5792),
            .I(visibleYZ0Z_2));
    Odrv4 I__1027 (
            .O(N__5789),
            .I(visibleYZ0Z_2));
    CascadeMux I__1026 (
            .O(N__5782),
            .I(N__5777));
    InMux I__1025 (
            .O(N__5781),
            .I(N__5774));
    InMux I__1024 (
            .O(N__5780),
            .I(N__5771));
    InMux I__1023 (
            .O(N__5777),
            .I(N__5768));
    LocalMux I__1022 (
            .O(N__5774),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0));
    LocalMux I__1021 (
            .O(N__5771),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0));
    LocalMux I__1020 (
            .O(N__5768),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0));
    InMux I__1019 (
            .O(N__5761),
            .I(N__5758));
    LocalMux I__1018 (
            .O(N__5758),
            .I(Pixel_RNOZ0Z_6));
    CascadeMux I__1017 (
            .O(N__5755),
            .I(un13_beamylt7_cascade_));
    InMux I__1016 (
            .O(N__5752),
            .I(N__5749));
    LocalMux I__1015 (
            .O(N__5749),
            .I(OutputEnabledZ0));
    InMux I__1014 (
            .O(N__5746),
            .I(N__5740));
    InMux I__1013 (
            .O(N__5745),
            .I(N__5740));
    LocalMux I__1012 (
            .O(N__5740),
            .I(N__5737));
    Odrv4 I__1011 (
            .O(N__5737),
            .I(un18_beamylt4));
    CascadeMux I__1010 (
            .O(N__5734),
            .I(un18_beamylto9_2_cascade_));
    InMux I__1009 (
            .O(N__5731),
            .I(N__5728));
    LocalMux I__1008 (
            .O(N__5728),
            .I(N__5725));
    Odrv4 I__1007 (
            .O(N__5725),
            .I(un8_beamy));
    CascadeMux I__1006 (
            .O(N__5722),
            .I(un18_beamylt10_0_cascade_));
    InMux I__1005 (
            .O(N__5719),
            .I(N__5716));
    LocalMux I__1004 (
            .O(N__5716),
            .I(N__5713));
    Odrv4 I__1003 (
            .O(N__5713),
            .I(un4_beamy_0));
    InMux I__1002 (
            .O(N__5710),
            .I(N__5707));
    LocalMux I__1001 (
            .O(N__5707),
            .I(un15_beamy_2));
    InMux I__1000 (
            .O(N__5704),
            .I(N__5701));
    LocalMux I__999 (
            .O(N__5701),
            .I(un13_beamylt7));
    CascadeMux I__998 (
            .O(N__5698),
            .I(un15_beamy_2_cascade_));
    IoInMux I__997 (
            .O(N__5695),
            .I(N__5692));
    LocalMux I__996 (
            .O(N__5692),
            .I(N__5689));
    Span4Mux_s2_h I__995 (
            .O(N__5689),
            .I(N__5686));
    Span4Mux_h I__994 (
            .O(N__5686),
            .I(N__5683));
    Odrv4 I__993 (
            .O(N__5683),
            .I(beamX_RNISO4TZ0Z_7));
    InMux I__992 (
            .O(N__5680),
            .I(N__5674));
    InMux I__991 (
            .O(N__5679),
            .I(N__5671));
    InMux I__990 (
            .O(N__5678),
            .I(N__5668));
    InMux I__989 (
            .O(N__5677),
            .I(N__5665));
    LocalMux I__988 (
            .O(N__5674),
            .I(beamYZ0Z_6));
    LocalMux I__987 (
            .O(N__5671),
            .I(beamYZ0Z_6));
    LocalMux I__986 (
            .O(N__5668),
            .I(beamYZ0Z_6));
    LocalMux I__985 (
            .O(N__5665),
            .I(beamYZ0Z_6));
    InMux I__984 (
            .O(N__5656),
            .I(N__5650));
    InMux I__983 (
            .O(N__5655),
            .I(N__5647));
    InMux I__982 (
            .O(N__5654),
            .I(N__5644));
    InMux I__981 (
            .O(N__5653),
            .I(N__5641));
    LocalMux I__980 (
            .O(N__5650),
            .I(beamYZ0Z_5));
    LocalMux I__979 (
            .O(N__5647),
            .I(beamYZ0Z_5));
    LocalMux I__978 (
            .O(N__5644),
            .I(beamYZ0Z_5));
    LocalMux I__977 (
            .O(N__5641),
            .I(beamYZ0Z_5));
    CascadeMux I__976 (
            .O(N__5632),
            .I(un4_beamylt6_cascade_));
    CascadeMux I__975 (
            .O(N__5629),
            .I(N__5624));
    InMux I__974 (
            .O(N__5628),
            .I(N__5619));
    InMux I__973 (
            .O(N__5627),
            .I(N__5616));
    InMux I__972 (
            .O(N__5624),
            .I(N__5611));
    InMux I__971 (
            .O(N__5623),
            .I(N__5611));
    InMux I__970 (
            .O(N__5622),
            .I(N__5608));
    LocalMux I__969 (
            .O(N__5619),
            .I(beamYZ0Z_9));
    LocalMux I__968 (
            .O(N__5616),
            .I(beamYZ0Z_9));
    LocalMux I__967 (
            .O(N__5611),
            .I(beamYZ0Z_9));
    LocalMux I__966 (
            .O(N__5608),
            .I(beamYZ0Z_9));
    InMux I__965 (
            .O(N__5599),
            .I(N__5592));
    InMux I__964 (
            .O(N__5598),
            .I(N__5589));
    InMux I__963 (
            .O(N__5597),
            .I(N__5584));
    InMux I__962 (
            .O(N__5596),
            .I(N__5584));
    InMux I__961 (
            .O(N__5595),
            .I(N__5581));
    LocalMux I__960 (
            .O(N__5592),
            .I(beamYZ0Z_8));
    LocalMux I__959 (
            .O(N__5589),
            .I(beamYZ0Z_8));
    LocalMux I__958 (
            .O(N__5584),
            .I(beamYZ0Z_8));
    LocalMux I__957 (
            .O(N__5581),
            .I(beamYZ0Z_8));
    CascadeMux I__956 (
            .O(N__5572),
            .I(un4_beamylt8_0_cascade_));
    InMux I__955 (
            .O(N__5569),
            .I(N__5561));
    InMux I__954 (
            .O(N__5568),
            .I(N__5558));
    InMux I__953 (
            .O(N__5567),
            .I(N__5555));
    InMux I__952 (
            .O(N__5566),
            .I(N__5550));
    InMux I__951 (
            .O(N__5565),
            .I(N__5550));
    InMux I__950 (
            .O(N__5564),
            .I(N__5547));
    LocalMux I__949 (
            .O(N__5561),
            .I(beamYZ0Z_7));
    LocalMux I__948 (
            .O(N__5558),
            .I(beamYZ0Z_7));
    LocalMux I__947 (
            .O(N__5555),
            .I(beamYZ0Z_7));
    LocalMux I__946 (
            .O(N__5550),
            .I(beamYZ0Z_7));
    LocalMux I__945 (
            .O(N__5547),
            .I(beamYZ0Z_7));
    InMux I__944 (
            .O(N__5536),
            .I(N__5529));
    InMux I__943 (
            .O(N__5535),
            .I(N__5523));
    InMux I__942 (
            .O(N__5534),
            .I(N__5518));
    InMux I__941 (
            .O(N__5533),
            .I(N__5518));
    InMux I__940 (
            .O(N__5532),
            .I(N__5515));
    LocalMux I__939 (
            .O(N__5529),
            .I(N__5512));
    InMux I__938 (
            .O(N__5528),
            .I(N__5507));
    InMux I__937 (
            .O(N__5527),
            .I(N__5507));
    InMux I__936 (
            .O(N__5526),
            .I(N__5504));
    LocalMux I__935 (
            .O(N__5523),
            .I(un5_vy));
    LocalMux I__934 (
            .O(N__5518),
            .I(un5_vy));
    LocalMux I__933 (
            .O(N__5515),
            .I(un5_vy));
    Odrv4 I__932 (
            .O(N__5512),
            .I(un5_vy));
    LocalMux I__931 (
            .O(N__5507),
            .I(un5_vy));
    LocalMux I__930 (
            .O(N__5504),
            .I(un5_vy));
    InMux I__929 (
            .O(N__5491),
            .I(N__5483));
    InMux I__928 (
            .O(N__5490),
            .I(N__5480));
    InMux I__927 (
            .O(N__5489),
            .I(N__5477));
    InMux I__926 (
            .O(N__5488),
            .I(N__5472));
    InMux I__925 (
            .O(N__5487),
            .I(N__5472));
    InMux I__924 (
            .O(N__5486),
            .I(N__5469));
    LocalMux I__923 (
            .O(N__5483),
            .I(beamYZ0Z_4));
    LocalMux I__922 (
            .O(N__5480),
            .I(beamYZ0Z_4));
    LocalMux I__921 (
            .O(N__5477),
            .I(beamYZ0Z_4));
    LocalMux I__920 (
            .O(N__5472),
            .I(beamYZ0Z_4));
    LocalMux I__919 (
            .O(N__5469),
            .I(beamYZ0Z_4));
    CascadeMux I__918 (
            .O(N__5458),
            .I(N__5455));
    InMux I__917 (
            .O(N__5455),
            .I(N__5452));
    LocalMux I__916 (
            .O(N__5452),
            .I(un8_beamylto9_1));
    CascadeMux I__915 (
            .O(N__5449),
            .I(N__5445));
    InMux I__914 (
            .O(N__5448),
            .I(N__5438));
    InMux I__913 (
            .O(N__5445),
            .I(N__5433));
    InMux I__912 (
            .O(N__5444),
            .I(N__5433));
    InMux I__911 (
            .O(N__5443),
            .I(N__5430));
    InMux I__910 (
            .O(N__5442),
            .I(N__5427));
    InMux I__909 (
            .O(N__5441),
            .I(N__5424));
    LocalMux I__908 (
            .O(N__5438),
            .I(beamYZ0Z_3));
    LocalMux I__907 (
            .O(N__5433),
            .I(beamYZ0Z_3));
    LocalMux I__906 (
            .O(N__5430),
            .I(beamYZ0Z_3));
    LocalMux I__905 (
            .O(N__5427),
            .I(beamYZ0Z_3));
    LocalMux I__904 (
            .O(N__5424),
            .I(beamYZ0Z_3));
    InMux I__903 (
            .O(N__5413),
            .I(N__5410));
    LocalMux I__902 (
            .O(N__5410),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41));
    CascadeMux I__901 (
            .O(N__5407),
            .I(Pixel_RNOZ0Z_5_cascade_));
    CascadeMux I__900 (
            .O(N__5404),
            .I(N_45_cascade_));
    InMux I__899 (
            .O(N__5401),
            .I(N__5398));
    LocalMux I__898 (
            .O(N__5398),
            .I(N_76));
    InMux I__897 (
            .O(N__5395),
            .I(N__5392));
    LocalMux I__896 (
            .O(N__5392),
            .I(TextOutputEnabledZ0));
    CascadeMux I__895 (
            .O(N__5389),
            .I(N_74_i_cascade_));
    IoInMux I__894 (
            .O(N__5386),
            .I(N__5383));
    LocalMux I__893 (
            .O(N__5383),
            .I(N__5380));
    IoSpan4Mux I__892 (
            .O(N__5380),
            .I(N__5377));
    Span4Mux_s2_v I__891 (
            .O(N__5377),
            .I(N__5374));
    Odrv4 I__890 (
            .O(N__5374),
            .I(Pixel_c));
    InMux I__889 (
            .O(N__5371),
            .I(N__5365));
    InMux I__888 (
            .O(N__5370),
            .I(N__5365));
    LocalMux I__887 (
            .O(N__5365),
            .I(N__5358));
    InMux I__886 (
            .O(N__5364),
            .I(N__5355));
    InMux I__885 (
            .O(N__5363),
            .I(N__5352));
    InMux I__884 (
            .O(N__5362),
            .I(N__5347));
    InMux I__883 (
            .O(N__5361),
            .I(N__5347));
    Odrv4 I__882 (
            .O(N__5358),
            .I(beamY_RNI9DLCZ0Z_2));
    LocalMux I__881 (
            .O(N__5355),
            .I(beamY_RNI9DLCZ0Z_2));
    LocalMux I__880 (
            .O(N__5352),
            .I(beamY_RNI9DLCZ0Z_2));
    LocalMux I__879 (
            .O(N__5347),
            .I(beamY_RNI9DLCZ0Z_2));
    CascadeMux I__878 (
            .O(N__5338),
            .I(N__5332));
    InMux I__877 (
            .O(N__5337),
            .I(N__5327));
    InMux I__876 (
            .O(N__5336),
            .I(N__5327));
    InMux I__875 (
            .O(N__5335),
            .I(N__5324));
    InMux I__874 (
            .O(N__5332),
            .I(N__5321));
    LocalMux I__873 (
            .O(N__5327),
            .I(beamYZ0Z_0));
    LocalMux I__872 (
            .O(N__5324),
            .I(beamYZ0Z_0));
    LocalMux I__871 (
            .O(N__5321),
            .I(beamYZ0Z_0));
    InMux I__870 (
            .O(N__5314),
            .I(N__5311));
    LocalMux I__869 (
            .O(N__5311),
            .I(un5_beamx_5));
    CascadeMux I__868 (
            .O(N__5308),
            .I(un1_beamy_4_cascade_));
    InMux I__867 (
            .O(N__5305),
            .I(N__5302));
    LocalMux I__866 (
            .O(N__5302),
            .I(un5_beamx_3));
    CascadeMux I__865 (
            .O(N__5299),
            .I(N__5296));
    InMux I__864 (
            .O(N__5296),
            .I(N__5289));
    InMux I__863 (
            .O(N__5295),
            .I(N__5284));
    InMux I__862 (
            .O(N__5294),
            .I(N__5284));
    InMux I__861 (
            .O(N__5293),
            .I(N__5279));
    InMux I__860 (
            .O(N__5292),
            .I(N__5279));
    LocalMux I__859 (
            .O(N__5289),
            .I(beamYZ0Z_1));
    LocalMux I__858 (
            .O(N__5284),
            .I(beamYZ0Z_1));
    LocalMux I__857 (
            .O(N__5279),
            .I(beamYZ0Z_1));
    CascadeMux I__856 (
            .O(N__5272),
            .I(N__5268));
    InMux I__855 (
            .O(N__5271),
            .I(N__5265));
    InMux I__854 (
            .O(N__5268),
            .I(N__5262));
    LocalMux I__853 (
            .O(N__5265),
            .I(un1_beamy_4));
    LocalMux I__852 (
            .O(N__5262),
            .I(un1_beamy_4));
    InMux I__851 (
            .O(N__5257),
            .I(N__5251));
    InMux I__850 (
            .O(N__5256),
            .I(N__5251));
    LocalMux I__849 (
            .O(N__5251),
            .I(un8_beamy_2));
    CascadeMux I__848 (
            .O(N__5248),
            .I(un1_beamylto9_2_cascade_));
    IoInMux I__847 (
            .O(N__5245),
            .I(N__5242));
    LocalMux I__846 (
            .O(N__5242),
            .I(N__5239));
    IoSpan4Mux I__845 (
            .O(N__5239),
            .I(N__5235));
    IoInMux I__844 (
            .O(N__5238),
            .I(N__5232));
    Sp12to4 I__843 (
            .O(N__5235),
            .I(N__5229));
    LocalMux I__842 (
            .O(N__5232),
            .I(N__5226));
    Span12Mux_v I__841 (
            .O(N__5229),
            .I(N__5223));
    Span4Mux_s2_v I__840 (
            .O(N__5226),
            .I(N__5220));
    Odrv12 I__839 (
            .O(N__5223),
            .I(VSync_c));
    Odrv4 I__838 (
            .O(N__5220),
            .I(VSync_c));
    InMux I__837 (
            .O(N__5215),
            .I(N__5212));
    LocalMux I__836 (
            .O(N__5212),
            .I(if_generate_plus_mult1_un68_sum_cry_2_s));
    InMux I__835 (
            .O(N__5209),
            .I(N__5203));
    InMux I__834 (
            .O(N__5208),
            .I(N__5203));
    LocalMux I__833 (
            .O(N__5203),
            .I(G_253));
    CascadeMux I__832 (
            .O(N__5200),
            .I(N__5197));
    InMux I__831 (
            .O(N__5197),
            .I(N__5194));
    LocalMux I__830 (
            .O(N__5194),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s));
    CascadeMux I__829 (
            .O(N__5191),
            .I(N__5186));
    InMux I__828 (
            .O(N__5190),
            .I(N__5182));
    InMux I__827 (
            .O(N__5189),
            .I(N__5175));
    InMux I__826 (
            .O(N__5186),
            .I(N__5175));
    InMux I__825 (
            .O(N__5185),
            .I(N__5175));
    LocalMux I__824 (
            .O(N__5182),
            .I(un9_r_0lto2));
    LocalMux I__823 (
            .O(N__5175),
            .I(un9_r_0lto2));
    InMux I__822 (
            .O(N__5170),
            .I(N__5167));
    LocalMux I__821 (
            .O(N__5167),
            .I(c_if_generate_plus_mult1_un75_sum_axbZ0Z_5));
    InMux I__820 (
            .O(N__5164),
            .I(c_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__819 (
            .O(N__5161),
            .I(N__5158));
    LocalMux I__818 (
            .O(N__5158),
            .I(N__5155));
    Odrv12 I__817 (
            .O(N__5155),
            .I(un9_r_1lt6_0));
    InMux I__816 (
            .O(N__5152),
            .I(N__5145));
    InMux I__815 (
            .O(N__5151),
            .I(N__5145));
    InMux I__814 (
            .O(N__5150),
            .I(N__5142));
    LocalMux I__813 (
            .O(N__5145),
            .I(N__5139));
    LocalMux I__812 (
            .O(N__5142),
            .I(N__5136));
    Span4Mux_v I__811 (
            .O(N__5139),
            .I(N__5133));
    Odrv4 I__810 (
            .O(N__5136),
            .I(c_if_generate_plus_mult1_un68_sum));
    Odrv4 I__809 (
            .O(N__5133),
            .I(c_if_generate_plus_mult1_un68_sum));
    CascadeMux I__808 (
            .O(N__5128),
            .I(N__5125));
    InMux I__807 (
            .O(N__5125),
            .I(N__5122));
    LocalMux I__806 (
            .O(N__5122),
            .I(c_if_generate_plus_mult1_un68_sum_iZ0));
    CascadeMux I__805 (
            .O(N__5119),
            .I(N__5115));
    InMux I__804 (
            .O(N__5118),
            .I(N__5111));
    InMux I__803 (
            .O(N__5115),
            .I(N__5107));
    InMux I__802 (
            .O(N__5114),
            .I(N__5104));
    LocalMux I__801 (
            .O(N__5111),
            .I(N__5101));
    InMux I__800 (
            .O(N__5110),
            .I(N__5098));
    LocalMux I__799 (
            .O(N__5107),
            .I(un9_r_0lto3));
    LocalMux I__798 (
            .O(N__5104),
            .I(un9_r_0lto3));
    Odrv4 I__797 (
            .O(N__5101),
            .I(un9_r_0lto3));
    LocalMux I__796 (
            .O(N__5098),
            .I(un9_r_0lto3));
    InMux I__795 (
            .O(N__5089),
            .I(N__5083));
    InMux I__794 (
            .O(N__5088),
            .I(N__5083));
    LocalMux I__793 (
            .O(N__5083),
            .I(un9_r_0lto3_i));
    CascadeMux I__792 (
            .O(N__5080),
            .I(N__5077));
    InMux I__791 (
            .O(N__5077),
            .I(N__5074));
    LocalMux I__790 (
            .O(N__5074),
            .I(N_404_i));
    InMux I__789 (
            .O(N__5071),
            .I(N__5065));
    InMux I__788 (
            .O(N__5070),
            .I(N__5065));
    LocalMux I__787 (
            .O(N__5065),
            .I(c_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__786 (
            .O(N__5062),
            .I(bfn_6_10_0_));
    InMux I__785 (
            .O(N__5059),
            .I(un5_vx_cry_8));
    CascadeMux I__784 (
            .O(N__5056),
            .I(CO3_0_cascade_));
    InMux I__783 (
            .O(N__5053),
            .I(N__5050));
    LocalMux I__782 (
            .O(N__5050),
            .I(N__5047));
    Span4Mux_h I__781 (
            .O(N__5047),
            .I(N__5044));
    Odrv4 I__780 (
            .O(N__5044),
            .I(N_14));
    CascadeMux I__779 (
            .O(N__5041),
            .I(N_3_0_cascade_));
    InMux I__778 (
            .O(N__5038),
            .I(N__5035));
    LocalMux I__777 (
            .O(N__5035),
            .I(N__5032));
    Odrv4 I__776 (
            .O(N__5032),
            .I(c_if_generate_plus_mult1_un75_sum));
    CascadeMux I__775 (
            .O(N__5029),
            .I(N__5024));
    CascadeMux I__774 (
            .O(N__5028),
            .I(N__5019));
    InMux I__773 (
            .O(N__5027),
            .I(N__5016));
    InMux I__772 (
            .O(N__5024),
            .I(N__5007));
    InMux I__771 (
            .O(N__5023),
            .I(N__5007));
    InMux I__770 (
            .O(N__5022),
            .I(N__5007));
    InMux I__769 (
            .O(N__5019),
            .I(N__5007));
    LocalMux I__768 (
            .O(N__5016),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0));
    LocalMux I__767 (
            .O(N__5007),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0));
    InMux I__766 (
            .O(N__5002),
            .I(un5_vx_cry_1));
    InMux I__765 (
            .O(N__4999),
            .I(un5_vx_cry_2));
    InMux I__764 (
            .O(N__4996),
            .I(N__4990));
    InMux I__763 (
            .O(N__4995),
            .I(N__4990));
    LocalMux I__762 (
            .O(N__4990),
            .I(N__4986));
    InMux I__761 (
            .O(N__4989),
            .I(N__4983));
    Span4Mux_h I__760 (
            .O(N__4986),
            .I(N__4980));
    LocalMux I__759 (
            .O(N__4983),
            .I(c_if_generate_plus_mult1_un61_sum));
    Odrv4 I__758 (
            .O(N__4980),
            .I(c_if_generate_plus_mult1_un61_sum));
    InMux I__757 (
            .O(N__4975),
            .I(un5_vx_cry_3));
    InMux I__756 (
            .O(N__4972),
            .I(un5_vx_cry_4));
    InMux I__755 (
            .O(N__4969),
            .I(un5_vx_cry_5));
    InMux I__754 (
            .O(N__4966),
            .I(un5_vx_cry_6));
    InMux I__753 (
            .O(N__4963),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6));
    CascadeMux I__752 (
            .O(N__4960),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41_cascade_));
    InMux I__751 (
            .O(N__4957),
            .I(N__4951));
    InMux I__750 (
            .O(N__4956),
            .I(N__4951));
    LocalMux I__749 (
            .O(N__4951),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7CZ0Z11));
    InMux I__748 (
            .O(N__4948),
            .I(N__4945));
    LocalMux I__747 (
            .O(N__4945),
            .I(Pixel_RNOZ0Z_7));
    InMux I__746 (
            .O(N__4942),
            .I(N__4938));
    InMux I__745 (
            .O(N__4941),
            .I(N__4935));
    LocalMux I__744 (
            .O(N__4938),
            .I(N__4930));
    LocalMux I__743 (
            .O(N__4935),
            .I(N__4930));
    Span4Mux_v I__742 (
            .O(N__4930),
            .I(N__4927));
    Odrv4 I__741 (
            .O(N__4927),
            .I(visibleYZ0Z_3));
    CascadeMux I__740 (
            .O(N__4924),
            .I(N__4921));
    InMux I__739 (
            .O(N__4921),
            .I(N__4918));
    LocalMux I__738 (
            .O(N__4918),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_0));
    CascadeMux I__737 (
            .O(N__4915),
            .I(N__4912));
    InMux I__736 (
            .O(N__4912),
            .I(N__4909));
    LocalMux I__735 (
            .O(N__4909),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000BZ0));
    InMux I__734 (
            .O(N__4906),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__733 (
            .O(N__4903),
            .I(N__4900));
    LocalMux I__732 (
            .O(N__4900),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73PZ0Z94));
    InMux I__731 (
            .O(N__4897),
            .I(N__4894));
    LocalMux I__730 (
            .O(N__4894),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SEZ0));
    InMux I__729 (
            .O(N__4891),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3));
    CascadeMux I__728 (
            .O(N__4888),
            .I(N__4884));
    InMux I__727 (
            .O(N__4887),
            .I(N__4875));
    InMux I__726 (
            .O(N__4884),
            .I(N__4875));
    InMux I__725 (
            .O(N__4883),
            .I(N__4875));
    InMux I__724 (
            .O(N__4882),
            .I(N__4872));
    LocalMux I__723 (
            .O(N__4875),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0));
    LocalMux I__722 (
            .O(N__4872),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0));
    CascadeMux I__721 (
            .O(N__4867),
            .I(N__4864));
    InMux I__720 (
            .O(N__4864),
            .I(N__4861));
    LocalMux I__719 (
            .O(N__4861),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQZ0Z56));
    InMux I__718 (
            .O(N__4858),
            .I(N__4855));
    LocalMux I__717 (
            .O(N__4855),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OGZ0));
    InMux I__716 (
            .O(N__4852),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__715 (
            .O(N__4849),
            .I(N__4846));
    LocalMux I__714 (
            .O(N__4846),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUTZ0Z97));
    CascadeMux I__713 (
            .O(N__4843),
            .I(N__4840));
    InMux I__712 (
            .O(N__4840),
            .I(N__4837));
    LocalMux I__711 (
            .O(N__4837),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_7));
    InMux I__710 (
            .O(N__4834),
            .I(N__4831));
    LocalMux I__709 (
            .O(N__4831),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_axb_7));
    InMux I__708 (
            .O(N__4828),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5));
    InMux I__707 (
            .O(N__4825),
            .I(N__4822));
    LocalMux I__706 (
            .O(N__4822),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_axb_7));
    InMux I__705 (
            .O(N__4819),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6));
    InMux I__704 (
            .O(N__4816),
            .I(un21_beamy_cry_8));
    InMux I__703 (
            .O(N__4813),
            .I(N__4810));
    LocalMux I__702 (
            .O(N__4810),
            .I(N__4807));
    Odrv4 I__701 (
            .O(N__4807),
            .I(if_generate_plus_mult1_un82_sum_s_5));
    CascadeMux I__700 (
            .O(N__4804),
            .I(N__4801));
    InMux I__699 (
            .O(N__4801),
            .I(N__4798));
    LocalMux I__698 (
            .O(N__4798),
            .I(un7_r_4));
    InMux I__697 (
            .O(N__4795),
            .I(N__4791));
    CascadeMux I__696 (
            .O(N__4794),
            .I(N__4787));
    LocalMux I__695 (
            .O(N__4791),
            .I(N__4783));
    InMux I__694 (
            .O(N__4790),
            .I(N__4780));
    InMux I__693 (
            .O(N__4787),
            .I(N__4775));
    InMux I__692 (
            .O(N__4786),
            .I(N__4775));
    Odrv4 I__691 (
            .O(N__4783),
            .I(if_generate_plus_mult1_un75_sum_s_5));
    LocalMux I__690 (
            .O(N__4780),
            .I(if_generate_plus_mult1_un75_sum_s_5));
    LocalMux I__689 (
            .O(N__4775),
            .I(if_generate_plus_mult1_un75_sum_s_5));
    InMux I__688 (
            .O(N__4768),
            .I(N__4765));
    LocalMux I__687 (
            .O(N__4765),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_0));
    InMux I__686 (
            .O(N__4762),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__685 (
            .O(N__4759),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__684 (
            .O(N__4756),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4));
    CascadeMux I__683 (
            .O(N__4753),
            .I(N__4750));
    InMux I__682 (
            .O(N__4750),
            .I(N__4747));
    LocalMux I__681 (
            .O(N__4747),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_7));
    InMux I__680 (
            .O(N__4744),
            .I(bfn_6_4_0_));
    InMux I__679 (
            .O(N__4741),
            .I(un21_beamy_cry_2));
    InMux I__678 (
            .O(N__4738),
            .I(un21_beamy_cry_3));
    InMux I__677 (
            .O(N__4735),
            .I(un21_beamy_cry_4));
    InMux I__676 (
            .O(N__4732),
            .I(un21_beamy_cry_5));
    InMux I__675 (
            .O(N__4729),
            .I(un21_beamy_cry_6));
    InMux I__674 (
            .O(N__4726),
            .I(un21_beamy_cry_7));
    CascadeMux I__673 (
            .O(N__4723),
            .I(N__4720));
    InMux I__672 (
            .O(N__4720),
            .I(N__4717));
    LocalMux I__671 (
            .O(N__4717),
            .I(if_generate_plus_mult1_un61_sum_cry_3_s));
    InMux I__670 (
            .O(N__4714),
            .I(c_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__669 (
            .O(N__4711),
            .I(N__4708));
    LocalMux I__668 (
            .O(N__4708),
            .I(c_if_generate_plus_mult1_un68_sum_axbZ0Z_5));
    InMux I__667 (
            .O(N__4705),
            .I(c_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__666 (
            .O(N__4702),
            .I(c_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__665 (
            .O(N__4699),
            .I(N__4693));
    InMux I__664 (
            .O(N__4698),
            .I(N__4693));
    LocalMux I__663 (
            .O(N__4693),
            .I(visibleYZ0Z_9));
    CascadeMux I__662 (
            .O(N__4690),
            .I(N__4687));
    InMux I__661 (
            .O(N__4687),
            .I(N__4684));
    LocalMux I__660 (
            .O(N__4684),
            .I(visibleY_RNIOR3DZ0Z_9));
    CascadeMux I__659 (
            .O(N__4681),
            .I(N__4678));
    InMux I__658 (
            .O(N__4678),
            .I(N__4675));
    LocalMux I__657 (
            .O(N__4675),
            .I(c_if_generate_plus_mult1_un61_sum_iZ0));
    InMux I__656 (
            .O(N__4672),
            .I(c_if_generate_plus_mult1_un68_sum_cry_1));
    InMux I__655 (
            .O(N__4669),
            .I(c_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__654 (
            .O(N__4666),
            .I(c_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__653 (
            .O(N__4663),
            .I(c_if_generate_plus_mult1_un68_sum_cry_4));
    CascadeMux I__652 (
            .O(N__4660),
            .I(N__4657));
    InMux I__651 (
            .O(N__4657),
            .I(N__4654));
    LocalMux I__650 (
            .O(N__4654),
            .I(if_generate_plus_mult1_un61_sum_cry_2_s));
    InMux I__649 (
            .O(N__4651),
            .I(c_if_generate_plus_mult1_un61_sum_cry_1));
    InMux I__648 (
            .O(N__4648),
            .I(N__4644));
    InMux I__647 (
            .O(N__4647),
            .I(N__4641));
    LocalMux I__646 (
            .O(N__4644),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32));
    LocalMux I__645 (
            .O(N__4641),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32));
    CascadeMux I__644 (
            .O(N__4636),
            .I(N__4633));
    InMux I__643 (
            .O(N__4633),
            .I(N__4630));
    LocalMux I__642 (
            .O(N__4630),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5KZ0Z3));
    InMux I__641 (
            .O(N__4627),
            .I(N__4624));
    LocalMux I__640 (
            .O(N__4624),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_axb_7));
    InMux I__639 (
            .O(N__4621),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5));
    InMux I__638 (
            .O(N__4618),
            .I(N__4615));
    LocalMux I__637 (
            .O(N__4615),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_axb_7));
    InMux I__636 (
            .O(N__4612),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6));
    CascadeMux I__635 (
            .O(N__4609),
            .I(N__4605));
    InMux I__634 (
            .O(N__4608),
            .I(N__4596));
    InMux I__633 (
            .O(N__4605),
            .I(N__4596));
    InMux I__632 (
            .O(N__4604),
            .I(N__4596));
    InMux I__631 (
            .O(N__4603),
            .I(N__4593));
    LocalMux I__630 (
            .O(N__4596),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3));
    LocalMux I__629 (
            .O(N__4593),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3));
    CascadeMux I__628 (
            .O(N__4588),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3_cascade_));
    CascadeMux I__627 (
            .O(N__4585),
            .I(N__4582));
    InMux I__626 (
            .O(N__4582),
            .I(N__4579));
    LocalMux I__625 (
            .O(N__4579),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_7));
    InMux I__624 (
            .O(N__4576),
            .I(N__4572));
    InMux I__623 (
            .O(N__4575),
            .I(N__4569));
    LocalMux I__622 (
            .O(N__4572),
            .I(visibleYZ0Z_8));
    LocalMux I__621 (
            .O(N__4569),
            .I(visibleYZ0Z_8));
    InMux I__620 (
            .O(N__4564),
            .I(N__4561));
    LocalMux I__619 (
            .O(N__4561),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJZ0));
    InMux I__618 (
            .O(N__4558),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2));
    InMux I__617 (
            .O(N__4555),
            .I(N__4552));
    LocalMux I__616 (
            .O(N__4552),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJZ0));
    InMux I__615 (
            .O(N__4549),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3));
    InMux I__614 (
            .O(N__4546),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5));
    InMux I__613 (
            .O(N__4543),
            .I(N__4540));
    LocalMux I__612 (
            .O(N__4540),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO));
    CascadeMux I__611 (
            .O(N__4537),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_));
    CascadeMux I__610 (
            .O(N__4534),
            .I(N__4529));
    CascadeMux I__609 (
            .O(N__4533),
            .I(N__4526));
    InMux I__608 (
            .O(N__4532),
            .I(N__4523));
    InMux I__607 (
            .O(N__4529),
            .I(N__4520));
    InMux I__606 (
            .O(N__4526),
            .I(N__4517));
    LocalMux I__605 (
            .O(N__4523),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__604 (
            .O(N__4520),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    LocalMux I__603 (
            .O(N__4517),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6));
    InMux I__602 (
            .O(N__4510),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5));
    InMux I__601 (
            .O(N__4507),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6));
    CascadeMux I__600 (
            .O(N__4504),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0_cascade_));
    InMux I__599 (
            .O(N__4501),
            .I(N__4495));
    InMux I__598 (
            .O(N__4500),
            .I(N__4495));
    LocalMux I__597 (
            .O(N__4495),
            .I(N__4492));
    Span4Mux_v I__596 (
            .O(N__4492),
            .I(N__4489));
    Odrv4 I__595 (
            .O(N__4489),
            .I(visibleYZ0Z_4));
    InMux I__594 (
            .O(N__4486),
            .I(N__4482));
    InMux I__593 (
            .O(N__4485),
            .I(N__4479));
    LocalMux I__592 (
            .O(N__4482),
            .I(N__4476));
    LocalMux I__591 (
            .O(N__4479),
            .I(N__4471));
    Span4Mux_v I__590 (
            .O(N__4476),
            .I(N__4471));
    Odrv4 I__589 (
            .O(N__4471),
            .I(visibleYZ0Z_5));
    CascadeMux I__588 (
            .O(N__4468),
            .I(N__4465));
    InMux I__587 (
            .O(N__4465),
            .I(N__4462));
    LocalMux I__586 (
            .O(N__4462),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_i_0));
    InMux I__585 (
            .O(N__4459),
            .I(N__4456));
    LocalMux I__584 (
            .O(N__4456),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSVZ0Z1));
    InMux I__583 (
            .O(N__4453),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__582 (
            .O(N__4450),
            .I(N__4447));
    LocalMux I__581 (
            .O(N__4447),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71EZ0Z1));
    CascadeMux I__580 (
            .O(N__4444),
            .I(N__4441));
    InMux I__579 (
            .O(N__4441),
            .I(N__4438));
    LocalMux I__578 (
            .O(N__4438),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0VZ0Z33));
    InMux I__577 (
            .O(N__4435),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3));
    CascadeMux I__576 (
            .O(N__4432),
            .I(N__4428));
    InMux I__575 (
            .O(N__4431),
            .I(N__4419));
    InMux I__574 (
            .O(N__4428),
            .I(N__4419));
    InMux I__573 (
            .O(N__4427),
            .I(N__4419));
    InMux I__572 (
            .O(N__4426),
            .I(N__4416));
    LocalMux I__571 (
            .O(N__4419),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1));
    LocalMux I__570 (
            .O(N__4416),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1));
    CascadeMux I__569 (
            .O(N__4411),
            .I(N__4408));
    InMux I__568 (
            .O(N__4408),
            .I(N__4405));
    LocalMux I__567 (
            .O(N__4405),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5TZ0Z1));
    InMux I__566 (
            .O(N__4402),
            .I(N__4399));
    LocalMux I__565 (
            .O(N__4399),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4JZ0Z3));
    InMux I__564 (
            .O(N__4396),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4));
    InMux I__563 (
            .O(N__4393),
            .I(N__4390));
    LocalMux I__562 (
            .O(N__4390),
            .I(un5_vy_cry_6_c_RNIG9KKZ0));
    InMux I__561 (
            .O(N__4387),
            .I(N__4384));
    LocalMux I__560 (
            .O(N__4384),
            .I(if_generate_plus_mult1_un47_sum_axb_4_l_ofx));
    InMux I__559 (
            .O(N__4381),
            .I(N__4378));
    LocalMux I__558 (
            .O(N__4378),
            .I(N__4372));
    InMux I__557 (
            .O(N__4377),
            .I(N__4365));
    InMux I__556 (
            .O(N__4376),
            .I(N__4365));
    InMux I__555 (
            .O(N__4375),
            .I(N__4365));
    Span4Mux_v I__554 (
            .O(N__4372),
            .I(N__4362));
    LocalMux I__553 (
            .O(N__4365),
            .I(N__4359));
    Odrv4 I__552 (
            .O(N__4362),
            .I(un5_vy_cry_6_c_RNI9MAAZ0));
    Odrv4 I__551 (
            .O(N__4359),
            .I(un5_vy_cry_6_c_RNI9MAAZ0));
    CascadeMux I__550 (
            .O(N__4354),
            .I(N__4351));
    InMux I__549 (
            .O(N__4351),
            .I(N__4348));
    LocalMux I__548 (
            .O(N__4348),
            .I(N_7_i));
    InMux I__547 (
            .O(N__4345),
            .I(N__4339));
    InMux I__546 (
            .O(N__4344),
            .I(N__4336));
    InMux I__545 (
            .O(N__4343),
            .I(N__4333));
    InMux I__544 (
            .O(N__4342),
            .I(N__4330));
    LocalMux I__543 (
            .O(N__4339),
            .I(if_generate_plus_mult1_un47_sum_s_5));
    LocalMux I__542 (
            .O(N__4336),
            .I(if_generate_plus_mult1_un47_sum_s_5));
    LocalMux I__541 (
            .O(N__4333),
            .I(if_generate_plus_mult1_un47_sum_s_5));
    LocalMux I__540 (
            .O(N__4330),
            .I(if_generate_plus_mult1_un47_sum_s_5));
    InMux I__539 (
            .O(N__4321),
            .I(N__4318));
    LocalMux I__538 (
            .O(N__4318),
            .I(r_if_generate_plus_mult1_un47_sum_i_5));
    InMux I__537 (
            .O(N__4315),
            .I(N__4312));
    LocalMux I__536 (
            .O(N__4312),
            .I(N__4307));
    CascadeMux I__535 (
            .O(N__4311),
            .I(N__4304));
    CascadeMux I__534 (
            .O(N__4310),
            .I(N__4301));
    Span4Mux_h I__533 (
            .O(N__4307),
            .I(N__4296));
    InMux I__532 (
            .O(N__4304),
            .I(N__4287));
    InMux I__531 (
            .O(N__4301),
            .I(N__4287));
    InMux I__530 (
            .O(N__4300),
            .I(N__4287));
    InMux I__529 (
            .O(N__4299),
            .I(N__4287));
    Span4Mux_v I__528 (
            .O(N__4296),
            .I(N__4282));
    LocalMux I__527 (
            .O(N__4287),
            .I(N__4282));
    Odrv4 I__526 (
            .O(N__4282),
            .I(un5_vy_cry_5_c_RNI7J9AZ0));
    CascadeMux I__525 (
            .O(N__4279),
            .I(N__4276));
    InMux I__524 (
            .O(N__4276),
            .I(N__4273));
    LocalMux I__523 (
            .O(N__4273),
            .I(un5_vy_i_24));
    CascadeMux I__522 (
            .O(N__4270),
            .I(N__4267));
    InMux I__521 (
            .O(N__4267),
            .I(N__4264));
    LocalMux I__520 (
            .O(N__4264),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__519 (
            .O(N__4261),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2));
    InMux I__518 (
            .O(N__4258),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__517 (
            .O(N__4255),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4));
    InMux I__516 (
            .O(N__4252),
            .I(un5_vy_cry_4));
    InMux I__515 (
            .O(N__4249),
            .I(un5_vy_cry_5));
    InMux I__514 (
            .O(N__4246),
            .I(un5_vy_cry_6));
    InMux I__513 (
            .O(N__4243),
            .I(N__4239));
    InMux I__512 (
            .O(N__4242),
            .I(N__4234));
    LocalMux I__511 (
            .O(N__4239),
            .I(N__4231));
    InMux I__510 (
            .O(N__4238),
            .I(N__4228));
    InMux I__509 (
            .O(N__4237),
            .I(N__4225));
    LocalMux I__508 (
            .O(N__4234),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    Odrv4 I__507 (
            .O(N__4231),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    LocalMux I__506 (
            .O(N__4228),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    LocalMux I__505 (
            .O(N__4225),
            .I(if_generate_plus_mult1_un61_sum_s_5));
    InMux I__504 (
            .O(N__4216),
            .I(N__4213));
    LocalMux I__503 (
            .O(N__4213),
            .I(N__4207));
    InMux I__502 (
            .O(N__4212),
            .I(N__4204));
    InMux I__501 (
            .O(N__4211),
            .I(N__4201));
    InMux I__500 (
            .O(N__4210),
            .I(N__4198));
    Odrv4 I__499 (
            .O(N__4207),
            .I(if_generate_plus_mult1_un68_sum_s_5));
    LocalMux I__498 (
            .O(N__4204),
            .I(if_generate_plus_mult1_un68_sum_s_5));
    LocalMux I__497 (
            .O(N__4201),
            .I(if_generate_plus_mult1_un68_sum_s_5));
    LocalMux I__496 (
            .O(N__4198),
            .I(if_generate_plus_mult1_un68_sum_s_5));
    InMux I__495 (
            .O(N__4189),
            .I(N__4182));
    InMux I__494 (
            .O(N__4188),
            .I(N__4182));
    InMux I__493 (
            .O(N__4187),
            .I(N__4179));
    LocalMux I__492 (
            .O(N__4182),
            .I(N__4176));
    LocalMux I__491 (
            .O(N__4179),
            .I(r_if_generate_plus_mult1_un54_sum));
    Odrv4 I__490 (
            .O(N__4176),
            .I(r_if_generate_plus_mult1_un54_sum));
    CascadeMux I__489 (
            .O(N__4171),
            .I(N__4168));
    InMux I__488 (
            .O(N__4168),
            .I(N__4165));
    LocalMux I__487 (
            .O(N__4165),
            .I(r_if_generate_plus_mult1_un54_sum_i_0));
    InMux I__486 (
            .O(N__4162),
            .I(N__4159));
    LocalMux I__485 (
            .O(N__4159),
            .I(r_if_generate_plus_mult1_un54_sum_i_5));
    InMux I__484 (
            .O(N__4156),
            .I(N__4150));
    InMux I__483 (
            .O(N__4155),
            .I(N__4147));
    InMux I__482 (
            .O(N__4154),
            .I(N__4144));
    InMux I__481 (
            .O(N__4153),
            .I(N__4141));
    LocalMux I__480 (
            .O(N__4150),
            .I(if_generate_plus_mult1_un54_sum_s_5_0));
    LocalMux I__479 (
            .O(N__4147),
            .I(if_generate_plus_mult1_un54_sum_s_5_0));
    LocalMux I__478 (
            .O(N__4144),
            .I(if_generate_plus_mult1_un54_sum_s_5_0));
    LocalMux I__477 (
            .O(N__4141),
            .I(if_generate_plus_mult1_un54_sum_s_5_0));
    CascadeMux I__476 (
            .O(N__4132),
            .I(N__4129));
    InMux I__475 (
            .O(N__4129),
            .I(N__4126));
    LocalMux I__474 (
            .O(N__4126),
            .I(un7_r_1));
    InMux I__473 (
            .O(N__4123),
            .I(N__4116));
    InMux I__472 (
            .O(N__4122),
            .I(N__4116));
    InMux I__471 (
            .O(N__4121),
            .I(N__4113));
    LocalMux I__470 (
            .O(N__4116),
            .I(N__4110));
    LocalMux I__469 (
            .O(N__4113),
            .I(N__4105));
    Span4Mux_h I__468 (
            .O(N__4110),
            .I(N__4105));
    Odrv4 I__467 (
            .O(N__4105),
            .I(r_if_generate_plus_mult1_un47_sum));
    CascadeMux I__466 (
            .O(N__4102),
            .I(N__4099));
    InMux I__465 (
            .O(N__4099),
            .I(N__4096));
    LocalMux I__464 (
            .O(N__4096),
            .I(r_if_generate_plus_mult1_un47_sum_i_0));
    CascadeMux I__463 (
            .O(N__4093),
            .I(N__4090));
    InMux I__462 (
            .O(N__4090),
            .I(N__4087));
    LocalMux I__461 (
            .O(N__4087),
            .I(r_if_generate_plus_mult1_un68_sum_i_0));
    CascadeMux I__460 (
            .O(N__4084),
            .I(N__4081));
    InMux I__459 (
            .O(N__4081),
            .I(N__4078));
    LocalMux I__458 (
            .O(N__4078),
            .I(if_generate_plus_mult1_un75_sum_cry_3_s));
    InMux I__457 (
            .O(N__4075),
            .I(r_if_generate_plus_mult1_un75_sum_cry_2));
    InMux I__456 (
            .O(N__4072),
            .I(N__4069));
    LocalMux I__455 (
            .O(N__4069),
            .I(r_if_generate_plus_mult1_un68_sum_i_5));
    CascadeMux I__454 (
            .O(N__4066),
            .I(N__4063));
    InMux I__453 (
            .O(N__4063),
            .I(N__4060));
    LocalMux I__452 (
            .O(N__4060),
            .I(if_generate_plus_mult1_un68_sum_cry_3_s_0));
    InMux I__451 (
            .O(N__4057),
            .I(N__4054));
    LocalMux I__450 (
            .O(N__4054),
            .I(r_if_generate_plus_mult1_un82_sum_axbZ0Z_5));
    InMux I__449 (
            .O(N__4051),
            .I(r_if_generate_plus_mult1_un75_sum_cry_3));
    InMux I__448 (
            .O(N__4048),
            .I(N__4045));
    LocalMux I__447 (
            .O(N__4045),
            .I(r_if_generate_plus_mult1_un75_sum_axbZ0Z_5));
    InMux I__446 (
            .O(N__4042),
            .I(r_if_generate_plus_mult1_un75_sum_cry_4));
    InMux I__445 (
            .O(N__4039),
            .I(N__4035));
    InMux I__444 (
            .O(N__4038),
            .I(N__4032));
    LocalMux I__443 (
            .O(N__4035),
            .I(N__4028));
    LocalMux I__442 (
            .O(N__4032),
            .I(N__4025));
    InMux I__441 (
            .O(N__4031),
            .I(N__4022));
    Odrv4 I__440 (
            .O(N__4028),
            .I(r_if_generate_plus_mult1_un75_sum));
    Odrv4 I__439 (
            .O(N__4025),
            .I(r_if_generate_plus_mult1_un75_sum));
    LocalMux I__438 (
            .O(N__4022),
            .I(r_if_generate_plus_mult1_un75_sum));
    InMux I__437 (
            .O(N__4015),
            .I(un5_vy_cry_0));
    InMux I__436 (
            .O(N__4012),
            .I(N__4009));
    LocalMux I__435 (
            .O(N__4009),
            .I(N__4004));
    InMux I__434 (
            .O(N__4008),
            .I(N__3999));
    InMux I__433 (
            .O(N__4007),
            .I(N__3999));
    Odrv4 I__432 (
            .O(N__4004),
            .I(r_if_generate_plus_mult1_un68_sum));
    LocalMux I__431 (
            .O(N__3999),
            .I(r_if_generate_plus_mult1_un68_sum));
    InMux I__430 (
            .O(N__3994),
            .I(un5_vy_cry_1));
    InMux I__429 (
            .O(N__3991),
            .I(N__3986));
    InMux I__428 (
            .O(N__3990),
            .I(N__3981));
    InMux I__427 (
            .O(N__3989),
            .I(N__3981));
    LocalMux I__426 (
            .O(N__3986),
            .I(r_if_generate_plus_mult1_un61_sum));
    LocalMux I__425 (
            .O(N__3981),
            .I(r_if_generate_plus_mult1_un61_sum));
    InMux I__424 (
            .O(N__3976),
            .I(un5_vy_cry_2));
    InMux I__423 (
            .O(N__3973),
            .I(un5_vy_cry_3));
    InMux I__422 (
            .O(N__3970),
            .I(N__3967));
    LocalMux I__421 (
            .O(N__3967),
            .I(visibleY_RNINQ3DZ0Z_8));
    InMux I__420 (
            .O(N__3964),
            .I(N__3961));
    LocalMux I__419 (
            .O(N__3961),
            .I(G_251));
    InMux I__418 (
            .O(N__3958),
            .I(N__3955));
    LocalMux I__417 (
            .O(N__3955),
            .I(G_252));
    InMux I__416 (
            .O(N__3952),
            .I(r_if_generate_plus_mult1_un82_sum_cry_4));
    InMux I__415 (
            .O(N__3949),
            .I(N__3943));
    InMux I__414 (
            .O(N__3948),
            .I(N__3943));
    LocalMux I__413 (
            .O(N__3943),
            .I(G_250));
    CascadeMux I__412 (
            .O(N__3940),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1_cascade_));
    InMux I__411 (
            .O(N__3937),
            .I(N__3933));
    InMux I__410 (
            .O(N__3936),
            .I(N__3930));
    LocalMux I__409 (
            .O(N__3933),
            .I(N__3927));
    LocalMux I__408 (
            .O(N__3930),
            .I(visibleYZ0Z_7));
    Odrv12 I__407 (
            .O(N__3927),
            .I(visibleYZ0Z_7));
    InMux I__406 (
            .O(N__3922),
            .I(N__3919));
    LocalMux I__405 (
            .O(N__3919),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450QZ0));
    InMux I__404 (
            .O(N__3916),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2));
    CascadeMux I__403 (
            .O(N__3913),
            .I(N__3910));
    InMux I__402 (
            .O(N__3910),
            .I(N__3907));
    LocalMux I__401 (
            .O(N__3907),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9MZ0Z01));
    InMux I__400 (
            .O(N__3904),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3));
    InMux I__399 (
            .O(N__3901),
            .I(N__3898));
    LocalMux I__398 (
            .O(N__3898),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDOZ0Z01));
    InMux I__397 (
            .O(N__3895),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4));
    InMux I__396 (
            .O(N__3892),
            .I(N__3889));
    LocalMux I__395 (
            .O(N__3889),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO));
    InMux I__394 (
            .O(N__3886),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5));
    InMux I__393 (
            .O(N__3883),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6));
    CascadeMux I__392 (
            .O(N__3880),
            .I(N__3875));
    InMux I__391 (
            .O(N__3879),
            .I(N__3865));
    InMux I__390 (
            .O(N__3878),
            .I(N__3865));
    InMux I__389 (
            .O(N__3875),
            .I(N__3865));
    InMux I__388 (
            .O(N__3874),
            .I(N__3865));
    LocalMux I__387 (
            .O(N__3865),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0));
    CascadeMux I__386 (
            .O(N__3862),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0_cascade_));
    CascadeMux I__385 (
            .O(N__3859),
            .I(N__3856));
    InMux I__384 (
            .O(N__3856),
            .I(N__3853));
    LocalMux I__383 (
            .O(N__3853),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_7));
    InMux I__382 (
            .O(N__3850),
            .I(r_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__381 (
            .O(N__3847),
            .I(N__3843));
    InMux I__380 (
            .O(N__3846),
            .I(N__3840));
    LocalMux I__379 (
            .O(N__3843),
            .I(N__3835));
    LocalMux I__378 (
            .O(N__3840),
            .I(N__3835));
    Odrv12 I__377 (
            .O(N__3835),
            .I(visibleYZ0Z_6));
    CascadeMux I__376 (
            .O(N__3832),
            .I(N__3829));
    InMux I__375 (
            .O(N__3829),
            .I(N__3826));
    LocalMux I__374 (
            .O(N__3826),
            .I(N__3823));
    Odrv4 I__373 (
            .O(N__3823),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_0));
    InMux I__372 (
            .O(N__3820),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__371 (
            .O(N__3817),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__370 (
            .O(N__3814),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4));
    InMux I__369 (
            .O(N__3811),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5));
    InMux I__368 (
            .O(N__3808),
            .I(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6));
    InMux I__367 (
            .O(N__3805),
            .I(N__3802));
    LocalMux I__366 (
            .O(N__3802),
            .I(N__3799));
    Odrv4 I__365 (
            .O(N__3799),
            .I(r_if_generate_plus_mult1_un68_sum_axbZ0Z_5));
    InMux I__364 (
            .O(N__3796),
            .I(r_if_generate_plus_mult1_un61_sum_cry_3));
    InMux I__363 (
            .O(N__3793),
            .I(r_if_generate_plus_mult1_un61_sum_cry_4));
    CascadeMux I__362 (
            .O(N__3790),
            .I(N__3787));
    InMux I__361 (
            .O(N__3787),
            .I(N__3784));
    LocalMux I__360 (
            .O(N__3784),
            .I(if_generate_plus_mult1_un54_sum_cry_3_s_0));
    InMux I__359 (
            .O(N__3781),
            .I(r_if_generate_plus_mult1_un54_sum_cry_2));
    InMux I__358 (
            .O(N__3778),
            .I(N__3775));
    LocalMux I__357 (
            .O(N__3775),
            .I(r_if_generate_plus_mult1_un61_sum_axbZ0Z_5));
    InMux I__356 (
            .O(N__3772),
            .I(r_if_generate_plus_mult1_un54_sum_cry_3));
    InMux I__355 (
            .O(N__3769),
            .I(r_if_generate_plus_mult1_un54_sum_cry_4));
    CascadeMux I__354 (
            .O(N__3766),
            .I(N__3763));
    InMux I__353 (
            .O(N__3763),
            .I(N__3760));
    LocalMux I__352 (
            .O(N__3760),
            .I(if_generate_plus_mult1_un47_sum_cry_3_s));
    InMux I__351 (
            .O(N__3757),
            .I(r_if_generate_plus_mult1_un47_sum_cry_2));
    InMux I__350 (
            .O(N__3754),
            .I(N__3751));
    LocalMux I__349 (
            .O(N__3751),
            .I(r_if_generate_plus_mult1_un54_sum_axbZ0Z_5));
    InMux I__348 (
            .O(N__3748),
            .I(r_if_generate_plus_mult1_un47_sum_cry_3));
    InMux I__347 (
            .O(N__3745),
            .I(r_if_generate_plus_mult1_un68_sum_cry_2));
    InMux I__346 (
            .O(N__3742),
            .I(r_if_generate_plus_mult1_un68_sum_cry_3));
    InMux I__345 (
            .O(N__3739),
            .I(r_if_generate_plus_mult1_un68_sum_cry_4));
    InMux I__344 (
            .O(N__3736),
            .I(N__3733));
    LocalMux I__343 (
            .O(N__3733),
            .I(r_if_generate_plus_mult1_un61_sum_i_5));
    CascadeMux I__342 (
            .O(N__3730),
            .I(N__3727));
    InMux I__341 (
            .O(N__3727),
            .I(N__3724));
    LocalMux I__340 (
            .O(N__3724),
            .I(r_if_generate_plus_mult1_un61_sum_i_0));
    CascadeMux I__339 (
            .O(N__3721),
            .I(N__3718));
    InMux I__338 (
            .O(N__3718),
            .I(N__3715));
    LocalMux I__337 (
            .O(N__3715),
            .I(N__3712));
    Odrv4 I__336 (
            .O(N__3712),
            .I(if_generate_plus_mult1_un61_sum_cry_3_s_0));
    InMux I__335 (
            .O(N__3709),
            .I(r_if_generate_plus_mult1_un61_sum_cry_2));
    IoInMux I__334 (
            .O(N__3706),
            .I(N__3703));
    LocalMux I__333 (
            .O(N__3703),
            .I(N__3700));
    Span4Mux_s1_h I__332 (
            .O(N__3700),
            .I(N__3697));
    Span4Mux_h I__331 (
            .O(N__3697),
            .I(N__3694));
    Span4Mux_v I__330 (
            .O(N__3694),
            .I(N__3691));
    Odrv4 I__329 (
            .O(N__3691),
            .I(\Clock50MHz.PixelClock ));
    IoInMux I__328 (
            .O(N__3688),
            .I(N__3685));
    LocalMux I__327 (
            .O(N__3685),
            .I(N__3682));
    IoSpan4Mux I__326 (
            .O(N__3682),
            .I(N__3679));
    Odrv4 I__325 (
            .O(N__3679),
            .I(Clock12MHz_c));
    INV INVPixelZ0C (
            .O(INVPixelZ0C_net),
            .I(N__7367));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(un8_beamx_cry_8),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(un5_vx_cry_7),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(un21_beamy_cry_1_THRU_CRY_6_THRU_CO),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_11_0_));
    ICE_GB \Clock50MHz.PLLOUTCORE_derived_clock_RNI49H9  (
            .USERSIGNALTOGLOBALBUFFER(N__3706),
            .GLOBALBUFFEROUTPUT(PixelClock_g));
    ICE_GB beamX_RNISO4T_0_7 (
            .USERSIGNALTOGLOBALBUFFER(N__5695),
            .GLOBALBUFFEROUTPUT(un15_beamy_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam visibleY_4_LC_4_3_0.C_ON=1'b1;
    defparam visibleY_4_LC_4_3_0.SEQ_MODE=4'b1000;
    defparam visibleY_4_LC_4_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_4_LC_4_3_0 (
            .in0(_gnd_net_),
            .in1(N__4007),
            .in2(_gnd_net_),
            .in3(N__4008),
            .lcout(visibleYZ0Z_4),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(r_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(N__7363),
            .ce(N__7295),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un68_sum_cry_3_s_LC_4_3_1.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un68_sum_cry_3_s_LC_4_3_1.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un68_sum_cry_3_s_LC_4_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_if_generate_plus_mult1_un68_sum_cry_3_s_LC_4_3_1 (
            .in0(_gnd_net_),
            .in1(N__4243),
            .in2(N__3730),
            .in3(N__3745),
            .lcout(if_generate_plus_mult1_un68_sum_cry_3_s_0),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(r_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un75_sum_axb_5_LC_4_3_2.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un75_sum_axb_5_LC_4_3_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un75_sum_axb_5_LC_4_3_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 r_if_generate_plus_mult1_un75_sum_axb_5_LC_4_3_2 (
            .in0(N__4211),
            .in1(N__3736),
            .in2(N__3721),
            .in3(N__3742),
            .lcout(r_if_generate_plus_mult1_un75_sum_axbZ0Z_5),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(r_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un68_sum_s_5_LC_4_3_3.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un68_sum_s_5_LC_4_3_3.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un68_sum_s_5_LC_4_3_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_if_generate_plus_mult1_un68_sum_s_5_LC_4_3_3 (
            .in0(_gnd_net_),
            .in1(N__3805),
            .in2(_gnd_net_),
            .in3(N__3739),
            .lcout(if_generate_plus_mult1_un68_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_4_4_2.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_4_4_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_4_4_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un61_sum_sbtinv_5_LC_4_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4237),
            .lcout(r_if_generate_plus_mult1_un61_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_5.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_5.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un61_sum_sbtinv_LC_4_4_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3991),
            .lcout(r_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un68_sum_sbtinv_5_LC_4_4_7.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un68_sum_sbtinv_5_LC_4_4_7.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un68_sum_sbtinv_5_LC_4_4_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un68_sum_sbtinv_5_LC_4_4_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4210),
            .lcout(r_if_generate_plus_mult1_un68_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_5_LC_4_5_0.C_ON=1'b1;
    defparam visibleY_5_LC_4_5_0.SEQ_MODE=4'b1000;
    defparam visibleY_5_LC_4_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_5_LC_4_5_0 (
            .in0(_gnd_net_),
            .in1(N__3989),
            .in2(_gnd_net_),
            .in3(N__3990),
            .lcout(visibleYZ0Z_5),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(r_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(N__7357),
            .ce(N__7292),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_5_1.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_5_1.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_5_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_if_generate_plus_mult1_un61_sum_cry_3_s_LC_4_5_1 (
            .in0(_gnd_net_),
            .in1(N__4155),
            .in2(N__4171),
            .in3(N__3709),
            .lcout(if_generate_plus_mult1_un61_sum_cry_3_s_0),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(r_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un68_sum_axb_5_LC_4_5_2.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un68_sum_axb_5_LC_4_5_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un68_sum_axb_5_LC_4_5_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 r_if_generate_plus_mult1_un68_sum_axb_5_LC_4_5_2 (
            .in0(N__4238),
            .in1(N__4162),
            .in2(N__3790),
            .in3(N__3796),
            .lcout(r_if_generate_plus_mult1_un68_sum_axbZ0Z_5),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(r_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un61_sum_s_5_LC_4_5_3.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un61_sum_s_5_LC_4_5_3.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un61_sum_s_5_LC_4_5_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_if_generate_plus_mult1_un61_sum_s_5_LC_4_5_3 (
            .in0(_gnd_net_),
            .in1(N__3778),
            .in2(_gnd_net_),
            .in3(N__3793),
            .lcout(if_generate_plus_mult1_un61_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_6_LC_4_6_0.C_ON=1'b1;
    defparam visibleY_6_LC_4_6_0.SEQ_MODE=4'b1000;
    defparam visibleY_6_LC_4_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_6_LC_4_6_0 (
            .in0(_gnd_net_),
            .in1(N__4188),
            .in2(_gnd_net_),
            .in3(N__4189),
            .lcout(visibleYZ0Z_6),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(r_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(N__7354),
            .ce(N__7289),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_6_1.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_6_1.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_6_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_6_1 (
            .in0(_gnd_net_),
            .in1(N__4344),
            .in2(N__4102),
            .in3(N__3781),
            .lcout(if_generate_plus_mult1_un54_sum_cry_3_s_0),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(r_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un61_sum_axb_5_LC_4_6_2.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un61_sum_axb_5_LC_4_6_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un61_sum_axb_5_LC_4_6_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 r_if_generate_plus_mult1_un61_sum_axb_5_LC_4_6_2 (
            .in0(N__4154),
            .in1(N__4321),
            .in2(N__3766),
            .in3(N__3772),
            .lcout(r_if_generate_plus_mult1_un61_sum_axbZ0Z_5),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(r_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un54_sum_s_5_LC_4_6_3.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un54_sum_s_5_LC_4_6_3.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un54_sum_s_5_LC_4_6_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_if_generate_plus_mult1_un54_sum_s_5_LC_4_6_3 (
            .in0(_gnd_net_),
            .in1(N__3754),
            .in2(_gnd_net_),
            .in3(N__3769),
            .lcout(if_generate_plus_mult1_un54_sum_s_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_7_LC_4_7_0.C_ON=1'b1;
    defparam visibleY_7_LC_4_7_0.SEQ_MODE=4'b1000;
    defparam visibleY_7_LC_4_7_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_7_LC_4_7_0 (
            .in0(_gnd_net_),
            .in1(N__4122),
            .in2(_gnd_net_),
            .in3(N__4123),
            .lcout(visibleYZ0Z_7),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(r_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(N__7353),
            .ce(N__7288),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_7_1.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_7_1 (
            .in0(_gnd_net_),
            .in1(N__4393),
            .in2(N__4279),
            .in3(N__3757),
            .lcout(if_generate_plus_mult1_un47_sum_cry_3_s),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(r_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un54_sum_axb_5_LC_4_7_2.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un54_sum_axb_5_LC_4_7_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un54_sum_axb_5_LC_4_7_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 r_if_generate_plus_mult1_un54_sum_axb_5_LC_4_7_2 (
            .in0(N__4343),
            .in1(N__4387),
            .in2(N__4354),
            .in3(N__3748),
            .lcout(r_if_generate_plus_mult1_un54_sum_axbZ0Z_5),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(r_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un47_sum_s_5_LC_4_7_3.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un47_sum_s_5_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un47_sum_s_5_LC_4_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un47_sum_s_5_LC_4_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3850),
            .lcout(if_generate_plus_mult1_un47_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_4_8_1.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_4_8_1.LUT_INIT=16'b0011001100110011;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_LC_4_8_1 (
            .in0(_gnd_net_),
            .in1(N__3936),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_4_8_3.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_4_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_4_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_sbtinv_LC_4_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3847),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0 (
            .in0(_gnd_net_),
            .in1(N__3846),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71E1_LC_4_9_1.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71E1_LC_4_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71E1_LC_4_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71E1_LC_4_9_1 (
            .in0(_gnd_net_),
            .in1(N__3874),
            .in2(N__3832),
            .in3(N__3820),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_sbtinv_RNIO71EZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_2),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5T1_LC_4_9_2.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5T1_LC_4_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5T1_LC_4_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5T1_LC_4_9_2 (
            .in0(_gnd_net_),
            .in1(N__3922),
            .in2(N__3880),
            .in3(N__3817),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3_c_RNIRT5TZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_3),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4T32_LC_4_9_3.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4T32_LC_4_9_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4T32_LC_4_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4T32_LC_4_9_3 (
            .in0(_gnd_net_),
            .in1(N__3878),
            .in2(N__3913),
            .in3(N__3814),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNID4TZ0Z32),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQP8K3_LC_4_9_4.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQP8K3_LC_4_9_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQP8K3_LC_4_9_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIQP8K3_LC_4_9_4 (
            .in0(N__4426),
            .in1(N__3901),
            .in2(N__3859),
            .in3(N__3811),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8G1_LC_4_9_5.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8G1_LC_4_9_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8G1_LC_4_9_5.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8G1_LC_4_9_5 (
            .in0(N__3892),
            .in1(N__3879),
            .in2(N__4534),
            .in3(N__3808),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1),
            .ltout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIAF8GZ0Z1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5K3_LC_4_9_6.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5K3_LC_4_9_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5K3_LC_4_9_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5K3_LC_4_9_6 (
            .in0(N__4648),
            .in1(_gnd_net_),
            .in2(N__3940),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNINJ5KZ0Z3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_4_10_0.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_4_10_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_4_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_LC_4_10_0 (
            .in0(_gnd_net_),
            .in1(N__3937),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450Q_LC_4_10_1.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450Q_LC_4_10_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450Q_LC_4_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450Q_LC_4_10_1 (
            .in0(_gnd_net_),
            .in1(N__3970),
            .in2(N__7779),
            .in3(N__3916),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2_c_RNI450QZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_2),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9M01_LC_4_10_2.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9M01_LC_4_10_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9M01_LC_4_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9M01_LC_4_10_2 (
            .in0(_gnd_net_),
            .in1(N__4564),
            .in2(N__7781),
            .in3(N__3904),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3_c_RNIL9MZ0Z01),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_3),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDO01_LC_4_10_3.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDO01_LC_4_10_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDO01_LC_4_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDO01_LC_4_10_3 (
            .in0(_gnd_net_),
            .in1(N__4555),
            .in2(N__7780),
            .in3(N__3895),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNINDOZ0Z01),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_4_10_4.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_4_10_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_4_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_LUT4_0_LC_4_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4533),
            .in3(N__3886),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_LC_4_10_5.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_LC_4_10_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_LC_4_10_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_LC_4_10_5 (
            .in0(_gnd_net_),
            .in1(N__4543),
            .in2(_gnd_net_),
            .in3(N__3883),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0),
            .ltout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_0_LC_4_10_6.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_0_LC_4_10_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_0_LC_4_10_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_RNI2ONJ_0_LC_4_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3862),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_RNINQ3D_8_LC_4_10_7.C_ON=1'b0;
    defparam visibleY_RNINQ3D_8_LC_4_10_7.SEQ_MODE=4'b0000;
    defparam visibleY_RNINQ3D_8_LC_4_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 visibleY_RNINQ3D_8_LC_4_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4576),
            .lcout(visibleY_RNINQ3DZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_8_LC_4_11_1.C_ON=1'b0;
    defparam visibleY_8_LC_4_11_1.SEQ_MODE=4'b1000;
    defparam visibleY_8_LC_4_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_8_LC_4_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4315),
            .lcout(visibleYZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7356),
            .ce(N__7287),
            .sr(_gnd_net_));
    defparam visibleY_9_LC_4_11_3.C_ON=1'b0;
    defparam visibleY_9_LC_4_11_3.SEQ_MODE=4'b1000;
    defparam visibleY_9_LC_4_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_9_LC_4_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4381),
            .lcout(visibleYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7356),
            .ce(N__7287),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_2_0.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_2_0.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_2_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 r_if_generate_plus_mult1_un82_sum_cry_2_c_LC_5_2_0 (
            .in0(_gnd_net_),
            .in1(N__3948),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(r_if_generate_plus_mult1_un82_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un82_sum_cry_3_c_inv_LC_5_2_1.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un82_sum_cry_3_c_inv_LC_5_2_1.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un82_sum_cry_3_c_inv_LC_5_2_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un82_sum_cry_3_c_inv_LC_5_2_1 (
            .in0(_gnd_net_),
            .in1(N__3964),
            .in2(N__4794),
            .in3(N__4038),
            .lcout(G_251),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un82_sum_cry_2),
            .carryout(r_if_generate_plus_mult1_un82_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_5_2_2.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_5_2_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_5_2_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un82_sum_cry_4_c_inv_LC_5_2_2 (
            .in0(_gnd_net_),
            .in1(N__3958),
            .in2(N__4084),
            .in3(N__4786),
            .lcout(G_252),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un82_sum_cry_3),
            .carryout(r_if_generate_plus_mult1_un82_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un82_sum_s_5_LC_5_2_3.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un82_sum_s_5_LC_5_2_3.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un82_sum_s_5_LC_5_2_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_if_generate_plus_mult1_un82_sum_s_5_LC_5_2_3 (
            .in0(_gnd_net_),
            .in1(N__4057),
            .in2(_gnd_net_),
            .in3(N__3952),
            .lcout(if_generate_plus_mult1_un82_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_5_2_6.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_5_2_6.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_5_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un82_sum_cry_2_c_inv_LC_5_2_6 (
            .in0(N__7706),
            .in1(N__3949),
            .in2(_gnd_net_),
            .in3(N__5536),
            .lcout(G_250),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un68_sum_sbtinv_LC_5_2_7.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un68_sum_sbtinv_LC_5_2_7.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un68_sum_sbtinv_LC_5_2_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un68_sum_sbtinv_LC_5_2_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4012),
            .lcout(r_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_3_LC_5_3_0.C_ON=1'b1;
    defparam visibleY_3_LC_5_3_0.SEQ_MODE=4'b1000;
    defparam visibleY_3_LC_5_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_3_LC_5_3_0 (
            .in0(_gnd_net_),
            .in1(N__4031),
            .in2(_gnd_net_),
            .in3(N__4039),
            .lcout(visibleYZ0Z_3),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(r_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(N__7369),
            .ce(N__7299),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_3_1.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_3_1.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_3_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 r_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_3_1 (
            .in0(_gnd_net_),
            .in1(N__4212),
            .in2(N__4093),
            .in3(N__4075),
            .lcout(if_generate_plus_mult1_un75_sum_cry_3_s),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(r_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un82_sum_axb_5_LC_5_3_2.C_ON=1'b1;
    defparam r_if_generate_plus_mult1_un82_sum_axb_5_LC_5_3_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un82_sum_axb_5_LC_5_3_2.LUT_INIT=16'b1001011001101001;
    LogicCell40 r_if_generate_plus_mult1_un82_sum_axb_5_LC_5_3_2 (
            .in0(N__4790),
            .in1(N__4072),
            .in2(N__4066),
            .in3(N__4051),
            .lcout(r_if_generate_plus_mult1_un82_sum_axbZ0Z_5),
            .ltout(),
            .carryin(r_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(r_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un75_sum_s_5_LC_5_3_3.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un75_sum_s_5_LC_5_3_3.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un75_sum_s_5_LC_5_3_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 r_if_generate_plus_mult1_un75_sum_s_5_LC_5_3_3 (
            .in0(_gnd_net_),
            .in1(N__4048),
            .in2(_gnd_net_),
            .in3(N__4042),
            .lcout(if_generate_plus_mult1_un75_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_0_c_LC_5_4_0.C_ON=1'b1;
    defparam un5_vy_cry_0_c_LC_5_4_0.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_0_c_LC_5_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_vy_cry_0_c_LC_5_4_0 (
            .in0(_gnd_net_),
            .in1(N__5526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(un5_vy_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_0_c_RNIT34A_LC_5_4_1.C_ON=1'b1;
    defparam un5_vy_cry_0_c_RNIT34A_LC_5_4_1.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_0_c_RNIT34A_LC_5_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_vy_cry_0_c_RNIT34A_LC_5_4_1 (
            .in0(_gnd_net_),
            .in1(N__5441),
            .in2(_gnd_net_),
            .in3(N__4015),
            .lcout(r_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_vy_cry_0),
            .carryout(un5_vy_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_1_c_RNIV65A_LC_5_4_2.C_ON=1'b1;
    defparam un5_vy_cry_1_c_RNIV65A_LC_5_4_2.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_1_c_RNIV65A_LC_5_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_vy_cry_1_c_RNIV65A_LC_5_4_2 (
            .in0(_gnd_net_),
            .in1(N__5486),
            .in2(_gnd_net_),
            .in3(N__3994),
            .lcout(r_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_vy_cry_1),
            .carryout(un5_vy_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_2_c_RNI1A6A_LC_5_4_3.C_ON=1'b1;
    defparam un5_vy_cry_2_c_RNI1A6A_LC_5_4_3.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_2_c_RNI1A6A_LC_5_4_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_vy_cry_2_c_RNI1A6A_LC_5_4_3 (
            .in0(_gnd_net_),
            .in1(N__5653),
            .in2(N__7702),
            .in3(N__3976),
            .lcout(r_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_vy_cry_2),
            .carryout(un5_vy_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_3_c_RNI3D7A_LC_5_4_4.C_ON=1'b1;
    defparam un5_vy_cry_3_c_RNI3D7A_LC_5_4_4.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_3_c_RNI3D7A_LC_5_4_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_vy_cry_3_c_RNI3D7A_LC_5_4_4 (
            .in0(_gnd_net_),
            .in1(N__5677),
            .in2(N__7704),
            .in3(N__3973),
            .lcout(r_if_generate_plus_mult1_un54_sum),
            .ltout(),
            .carryin(un5_vy_cry_3),
            .carryout(un5_vy_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_4_c_RNI5G8A_LC_5_4_5.C_ON=1'b1;
    defparam un5_vy_cry_4_c_RNI5G8A_LC_5_4_5.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_4_c_RNI5G8A_LC_5_4_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_vy_cry_4_c_RNI5G8A_LC_5_4_5 (
            .in0(_gnd_net_),
            .in1(N__5564),
            .in2(N__7703),
            .in3(N__4252),
            .lcout(r_if_generate_plus_mult1_un47_sum),
            .ltout(),
            .carryin(un5_vy_cry_4),
            .carryout(un5_vy_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_5_c_RNI7J9A_LC_5_4_6.C_ON=1'b1;
    defparam un5_vy_cry_5_c_RNI7J9A_LC_5_4_6.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_5_c_RNI7J9A_LC_5_4_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_vy_cry_5_c_RNI7J9A_LC_5_4_6 (
            .in0(_gnd_net_),
            .in1(N__5595),
            .in2(N__7705),
            .in3(N__4249),
            .lcout(un5_vy_cry_5_c_RNI7J9AZ0),
            .ltout(),
            .carryin(un5_vy_cry_5),
            .carryout(un5_vy_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_6_c_RNI9MAA_LC_5_4_7.C_ON=1'b0;
    defparam un5_vy_cry_6_c_RNI9MAA_LC_5_4_7.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_6_c_RNI9MAA_LC_5_4_7.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_vy_cry_6_c_RNI9MAA_LC_5_4_7 (
            .in0(_gnd_net_),
            .in1(N__5622),
            .in2(_gnd_net_),
            .in3(N__4246),
            .lcout(un5_vy_cry_6_c_RNI9MAAZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TextOutputEnabled_RNO_0_LC_5_5_1.C_ON=1'b0;
    defparam TextOutputEnabled_RNO_0_LC_5_5_1.SEQ_MODE=4'b0000;
    defparam TextOutputEnabled_RNO_0_LC_5_5_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 TextOutputEnabled_RNO_0_LC_5_5_1 (
            .in0(N__6085),
            .in1(N__4242),
            .in2(N__4132),
            .in3(N__4216),
            .lcout(un7_r_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_5_2.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_5_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_5_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4187),
            .lcout(r_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_5_7.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_5_7.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_5_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_5_5_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4153),
            .lcout(r_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TextOutputEnabled_RNO_2_LC_5_6_5.C_ON=1'b0;
    defparam TextOutputEnabled_RNO_2_LC_5_6_5.SEQ_MODE=4'b0000;
    defparam TextOutputEnabled_RNO_2_LC_5_6_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 TextOutputEnabled_RNO_2_LC_5_6_5 (
            .in0(N__5053),
            .in1(N__4156),
            .in2(_gnd_net_),
            .in3(N__4345),
            .lcout(un7_r_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un47_sum_sbtinv_LC_5_6_6.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un47_sum_sbtinv_LC_5_6_6.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un47_sum_sbtinv_LC_5_6_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un47_sum_sbtinv_LC_5_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4121),
            .lcout(r_if_generate_plus_mult1_un47_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_7_0.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_7_0.LUT_INIT=16'b0011001100110011;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_LC_5_7_0 (
            .in0(_gnd_net_),
            .in1(N__4485),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_6_c_RNIG9KK_LC_5_7_1.C_ON=1'b0;
    defparam un5_vy_cry_6_c_RNIG9KK_LC_5_7_1.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_6_c_RNIG9KK_LC_5_7_1.LUT_INIT=16'b0011001111111111;
    LogicCell40 un5_vy_cry_6_c_RNIG9KK_LC_5_7_1 (
            .in0(_gnd_net_),
            .in1(N__4300),
            .in2(_gnd_net_),
            .in3(N__4375),
            .lcout(un5_vy_cry_6_c_RNIG9KKZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un47_sum_axb_4_l_ofx_LC_5_7_2.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un47_sum_axb_4_l_ofx_LC_5_7_2.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un47_sum_axb_4_l_ofx_LC_5_7_2.LUT_INIT=16'b1010000010100000;
    LogicCell40 r_if_generate_plus_mult1_un47_sum_axb_4_l_ofx_LC_5_7_2 (
            .in0(N__4376),
            .in1(_gnd_net_),
            .in2(N__4310),
            .in3(_gnd_net_),
            .lcout(if_generate_plus_mult1_un47_sum_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_6_c_RNIG9KK_0_LC_5_7_4.C_ON=1'b0;
    defparam un5_vy_cry_6_c_RNIG9KK_0_LC_5_7_4.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_6_c_RNIG9KK_0_LC_5_7_4.LUT_INIT=16'b0101101001011010;
    LogicCell40 un5_vy_cry_6_c_RNIG9KK_0_LC_5_7_4 (
            .in0(N__4377),
            .in1(_gnd_net_),
            .in2(N__4311),
            .in3(_gnd_net_),
            .lcout(N_7_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_if_generate_plus_mult1_un47_sum_sbtinv_5_LC_5_7_5.C_ON=1'b0;
    defparam r_if_generate_plus_mult1_un47_sum_sbtinv_5_LC_5_7_5.SEQ_MODE=4'b0000;
    defparam r_if_generate_plus_mult1_un47_sum_sbtinv_5_LC_5_7_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 r_if_generate_plus_mult1_un47_sum_sbtinv_5_LC_5_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4342),
            .lcout(r_if_generate_plus_mult1_un47_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vy_cry_5_c_RNI7J9A_0_LC_5_7_7.C_ON=1'b0;
    defparam un5_vy_cry_5_c_RNI7J9A_0_LC_5_7_7.SEQ_MODE=4'b0000;
    defparam un5_vy_cry_5_c_RNI7J9A_0_LC_5_7_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_vy_cry_5_c_RNI7J9A_0_LC_5_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4299),
            .lcout(un5_vy_i_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0 (
            .in0(_gnd_net_),
            .in1(N__4500),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73P94_LC_5_8_1.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73P94_LC_5_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73P94_LC_5_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73P94_LC_5_8_1 (
            .in0(_gnd_net_),
            .in1(N__4604),
            .in2(N__4270),
            .in3(N__4261),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_sbtinv_RNI73PZ0Z94),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQ56_LC_5_8_2.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQ56_LC_5_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQ56_LC_5_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQ56_LC_5_8_2 (
            .in0(_gnd_net_),
            .in1(N__4459),
            .in2(N__4609),
            .in3(N__4258),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3_c_RNI6HQZ0Z56),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUT97_LC_5_8_3.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUT97_LC_5_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUT97_LC_5_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUT97_LC_5_8_3 (
            .in0(_gnd_net_),
            .in1(N__4608),
            .in2(N__4444),
            .in3(N__4255),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNINUTZ0Z97),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIP00TH_LC_5_8_4.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIP00TH_LC_5_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIP00TH_LC_5_8_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIP00TH_LC_5_8_4 (
            .in0(N__4882),
            .in1(N__4402),
            .in2(N__4585),
            .in3(N__4510),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_LC_5_8_5.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_LC_5_8_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_LC_5_8_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_LC_5_8_5 (
            .in0(_gnd_net_),
            .in1(N__4627),
            .in2(_gnd_net_),
            .in3(N__4507),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0),
            .ltout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3AZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_0_LC_5_8_6.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_0_LC_5_8_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_0_LC_5_8_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNIT7R3A_0_LC_5_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4504),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_5_8_7.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_5_8_7.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_5_8_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_LC_5_8_7 (
            .in0(N__4501),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_9_0.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_9_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_LC_5_9_0 (
            .in0(_gnd_net_),
            .in1(N__4486),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSV1_LC_5_9_1.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSV1_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSV1_LC_5_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSV1_LC_5_9_1 (
            .in0(_gnd_net_),
            .in1(N__4427),
            .in2(N__4468),
            .in3(N__4453),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2_c_RNI5LSVZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0V33_LC_5_9_2.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0V33_LC_5_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0V33_LC_5_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0V33_LC_5_9_2 (
            .in0(_gnd_net_),
            .in1(N__4450),
            .in2(N__4432),
            .in3(N__4435),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3_c_RNIL0VZ0Z33),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4J3_LC_5_9_3.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4J3_LC_5_9_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4J3_LC_5_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4J3_LC_5_9_3 (
            .in0(_gnd_net_),
            .in1(N__4431),
            .in2(N__4411),
            .in3(N__4396),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNIPO4JZ0Z3),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI9FRN9_LC_5_9_4.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI9FRN9_LC_5_9_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI9FRN9_LC_5_9_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNI9FRN9_LC_5_9_4 (
            .in0(N__4603),
            .in1(N__4647),
            .in2(N__4636),
            .in3(N__4621),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_LC_5_9_5.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_LC_5_9_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_LC_5_9_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_LC_5_9_5 (
            .in0(_gnd_net_),
            .in1(N__4618),
            .in2(_gnd_net_),
            .in3(N__4612),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3),
            .ltout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91QZ0Z3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_0_LC_5_9_6.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_0_LC_5_9_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_0_LC_5_9_6.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNIG91Q3_0_LC_5_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4588),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un54_sum_i_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_5_10_0.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_5_10_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_5_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_LC_5_10_0 (
            .in0(_gnd_net_),
            .in1(N__4575),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJ_LC_5_10_1.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJ_LC_5_10_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJ_LC_5_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJ_LC_5_10_1 (
            .in0(_gnd_net_),
            .in1(N__7753),
            .in2(N__4690),
            .in3(N__4558),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2_c_RNI7TOJZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_2),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJ_LC_5_10_2.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJ_LC_5_10_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJ_LC_5_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJ_LC_5_10_2 (
            .in0(_gnd_net_),
            .in1(N__4699),
            .in2(N__7778),
            .in3(N__4549),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3_c_RNI8VPJZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_3),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_5_10_3.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_5_10_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_5_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_LUT4_0_LC_5_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4546),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO),
            .ltout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un33_sum_cry_5_THRU_CO_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_5_10_4.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_5_10_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_5_10_4.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_cry_6_c_inv_LC_5_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4537),
            .in3(N__4532),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un40_sum_axb_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_RNIOR3D_9_LC_5_10_6.C_ON=1'b0;
    defparam visibleY_RNIOR3D_9_LC_5_10_6.SEQ_MODE=4'b0000;
    defparam visibleY_RNIOR3D_9_LC_5_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 visibleY_RNIOR3D_9_LC_5_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4698),
            .lcout(visibleY_RNIOR3DZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un61_sum_i_LC_5_10_7.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un61_sum_i_LC_5_10_7.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un61_sum_i_LC_5_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 c_if_generate_plus_mult1_un61_sum_i_LC_5_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4989),
            .lcout(c_if_generate_plus_mult1_un61_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_3_LC_5_11_0.C_ON=1'b1;
    defparam visibleX_3_LC_5_11_0.SEQ_MODE=4'b1000;
    defparam visibleX_3_LC_5_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleX_3_LC_5_11_0 (
            .in0(_gnd_net_),
            .in1(N__5151),
            .in2(_gnd_net_),
            .in3(N__5152),
            .lcout(N_84),
            .ltout(),
            .carryin(bfn_5_11_0_),
            .carryout(c_if_generate_plus_mult1_un68_sum_cry_1),
            .clk(N__7359),
            .ce(N__7290),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un68_sum_cry_2_s_LC_5_11_1.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un68_sum_cry_2_s_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un68_sum_cry_2_s_LC_5_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un68_sum_cry_2_s_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(N__5088),
            .in2(N__4681),
            .in3(N__4672),
            .lcout(if_generate_plus_mult1_un68_sum_cry_2_s),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un68_sum_cry_1),
            .carryout(c_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_11_2.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_11_2.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_11_2 (
            .in0(_gnd_net_),
            .in1(N__5114),
            .in2(N__4660),
            .in3(N__4669),
            .lcout(if_generate_plus_mult1_un68_sum_cry_3_s),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(c_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un75_sum_axb_5_LC_5_11_3.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un75_sum_axb_5_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un75_sum_axb_5_LC_5_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 c_if_generate_plus_mult1_un75_sum_axb_5_LC_5_11_3 (
            .in0(N__5190),
            .in1(N__5089),
            .in2(N__4723),
            .in3(N__4666),
            .lcout(c_if_generate_plus_mult1_un75_sum_axbZ0Z_5),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(c_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un68_sum_s_5_LC_5_11_4.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un68_sum_s_5_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un68_sum_s_5_LC_5_11_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 c_if_generate_plus_mult1_un68_sum_s_5_LC_5_11_4 (
            .in0(_gnd_net_),
            .in1(N__4711),
            .in2(_gnd_net_),
            .in3(N__4663),
            .lcout(un9_r_0lto2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_4_LC_5_12_0.C_ON=1'b1;
    defparam visibleX_4_LC_5_12_0.SEQ_MODE=4'b1000;
    defparam visibleX_4_LC_5_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleX_4_LC_5_12_0 (
            .in0(_gnd_net_),
            .in1(N__4995),
            .in2(_gnd_net_),
            .in3(N__4996),
            .lcout(visibleXZ0Z_4),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(c_if_generate_plus_mult1_un61_sum_cry_1),
            .clk(N__7364),
            .ce(N__7293),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_12_1.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un61_sum_cry_2_s_LC_5_12_1 (
            .in0(_gnd_net_),
            .in1(N__5070),
            .in2(N__5080),
            .in3(N__4651),
            .lcout(if_generate_plus_mult1_un61_sum_cry_2_s),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un61_sum_cry_1),
            .carryout(c_if_generate_plus_mult1_un61_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_12_2.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_12_2 (
            .in0(_gnd_net_),
            .in1(N__6078),
            .in2(N__6196),
            .in3(N__4714),
            .lcout(if_generate_plus_mult1_un61_sum_cry_3_s),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un61_sum_cry_2),
            .carryout(c_if_generate_plus_mult1_un61_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un68_sum_axb_5_LC_5_12_3.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un68_sum_axb_5_LC_5_12_3.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un68_sum_axb_5_LC_5_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 c_if_generate_plus_mult1_un68_sum_axb_5_LC_5_12_3 (
            .in0(N__5118),
            .in1(N__5071),
            .in2(N__6157),
            .in3(N__4705),
            .lcout(c_if_generate_plus_mult1_un68_sum_axbZ0Z_5),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un61_sum_cry_3),
            .carryout(c_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un61_sum_s_5_LC_5_12_4.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un61_sum_s_5_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un61_sum_s_5_LC_5_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 c_if_generate_plus_mult1_un61_sum_s_5_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(N__6106),
            .in2(_gnd_net_),
            .in3(N__4702),
            .lcout(un9_r_0lto3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleY_1_LC_6_3_0.C_ON=1'b1;
    defparam visibleY_1_LC_6_3_0.SEQ_MODE=4'b1000;
    defparam visibleY_1_LC_6_3_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleY_1_LC_6_3_0 (
            .in0(_gnd_net_),
            .in1(N__5292),
            .in2(N__5338),
            .in3(N__5293),
            .lcout(visibleYZ0Z_1),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(un21_beamy_cry_1),
            .clk(N__7371),
            .ce(N__7300),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_THRU_CRY_0_LC_6_3_1.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_THRU_CRY_0_LC_6_3_1.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_THRU_CRY_0_LC_6_3_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_THRU_CRY_0_LC_6_3_1 (
            .in0(_gnd_net_),
            .in1(N__7723),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un21_beamy_cry_1),
            .carryout(un21_beamy_cry_1_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_THRU_CRY_1_LC_6_3_2.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_THRU_CRY_1_LC_6_3_2.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_THRU_CRY_1_LC_6_3_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_THRU_CRY_1_LC_6_3_2 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__7766),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un21_beamy_cry_1_THRU_CRY_0_THRU_CO),
            .carryout(un21_beamy_cry_1_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_THRU_CRY_2_LC_6_3_3.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_THRU_CRY_2_LC_6_3_3.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_THRU_CRY_2_LC_6_3_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_THRU_CRY_2_LC_6_3_3 (
            .in0(_gnd_net_),
            .in1(N__7727),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un21_beamy_cry_1_THRU_CRY_1_THRU_CO),
            .carryout(un21_beamy_cry_1_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_THRU_CRY_3_LC_6_3_4.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_THRU_CRY_3_LC_6_3_4.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_THRU_CRY_3_LC_6_3_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_THRU_CRY_3_LC_6_3_4 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__7767),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un21_beamy_cry_1_THRU_CRY_2_THRU_CO),
            .carryout(un21_beamy_cry_1_THRU_CRY_3_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_THRU_CRY_4_LC_6_3_5.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_THRU_CRY_4_LC_6_3_5.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_THRU_CRY_4_LC_6_3_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_THRU_CRY_4_LC_6_3_5 (
            .in0(_gnd_net_),
            .in1(N__7731),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un21_beamy_cry_1_THRU_CRY_3_THRU_CO),
            .carryout(un21_beamy_cry_1_THRU_CRY_4_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_THRU_CRY_5_LC_6_3_6.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_THRU_CRY_5_LC_6_3_6.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_THRU_CRY_5_LC_6_3_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_THRU_CRY_5_LC_6_3_6 (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__7768),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un21_beamy_cry_1_THRU_CRY_4_THRU_CO),
            .carryout(un21_beamy_cry_1_THRU_CRY_5_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un21_beamy_cry_1_c_THRU_CRY_6_LC_6_3_7.C_ON=1'b1;
    defparam un21_beamy_cry_1_c_THRU_CRY_6_LC_6_3_7.SEQ_MODE=4'b0000;
    defparam un21_beamy_cry_1_c_THRU_CRY_6_LC_6_3_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un21_beamy_cry_1_c_THRU_CRY_6_LC_6_3_7 (
            .in0(_gnd_net_),
            .in1(N__7735),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un21_beamy_cry_1_THRU_CRY_5_THRU_CO),
            .carryout(un21_beamy_cry_1_THRU_CRY_6_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_2_LC_6_4_0.C_ON=1'b1;
    defparam beamY_2_LC_6_4_0.SEQ_MODE=4'b1000;
    defparam beamY_2_LC_6_4_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_2_LC_6_4_0 (
            .in0(_gnd_net_),
            .in1(N__5532),
            .in2(_gnd_net_),
            .in3(N__4744),
            .lcout(un5_vy),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(un21_beamy_cry_2),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam beamY_3_LC_6_4_1.C_ON=1'b1;
    defparam beamY_3_LC_6_4_1.SEQ_MODE=4'b1000;
    defparam beamY_3_LC_6_4_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_3_LC_6_4_1 (
            .in0(N__5370),
            .in1(N__5448),
            .in2(_gnd_net_),
            .in3(N__4741),
            .lcout(beamYZ0Z_3),
            .ltout(),
            .carryin(un21_beamy_cry_2),
            .carryout(un21_beamy_cry_3),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam beamY_4_LC_6_4_2.C_ON=1'b1;
    defparam beamY_4_LC_6_4_2.SEQ_MODE=4'b1000;
    defparam beamY_4_LC_6_4_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_4_LC_6_4_2 (
            .in0(N__5361),
            .in1(N__5490),
            .in2(_gnd_net_),
            .in3(N__4738),
            .lcout(beamYZ0Z_4),
            .ltout(),
            .carryin(un21_beamy_cry_3),
            .carryout(un21_beamy_cry_4),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam beamY_5_LC_6_4_3.C_ON=1'b1;
    defparam beamY_5_LC_6_4_3.SEQ_MODE=4'b1000;
    defparam beamY_5_LC_6_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_5_LC_6_4_3 (
            .in0(_gnd_net_),
            .in1(N__5656),
            .in2(_gnd_net_),
            .in3(N__4735),
            .lcout(beamYZ0Z_5),
            .ltout(),
            .carryin(un21_beamy_cry_4),
            .carryout(un21_beamy_cry_5),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam beamY_6_LC_6_4_4.C_ON=1'b1;
    defparam beamY_6_LC_6_4_4.SEQ_MODE=4'b1000;
    defparam beamY_6_LC_6_4_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_6_LC_6_4_4 (
            .in0(_gnd_net_),
            .in1(N__5680),
            .in2(_gnd_net_),
            .in3(N__4732),
            .lcout(beamYZ0Z_6),
            .ltout(),
            .carryin(un21_beamy_cry_5),
            .carryout(un21_beamy_cry_6),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam beamY_7_LC_6_4_5.C_ON=1'b1;
    defparam beamY_7_LC_6_4_5.SEQ_MODE=4'b1000;
    defparam beamY_7_LC_6_4_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamY_7_LC_6_4_5 (
            .in0(N__5371),
            .in1(N__5568),
            .in2(_gnd_net_),
            .in3(N__4729),
            .lcout(beamYZ0Z_7),
            .ltout(),
            .carryin(un21_beamy_cry_6),
            .carryout(un21_beamy_cry_7),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam beamY_8_LC_6_4_6.C_ON=1'b1;
    defparam beamY_8_LC_6_4_6.SEQ_MODE=4'b1000;
    defparam beamY_8_LC_6_4_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamY_8_LC_6_4_6 (
            .in0(_gnd_net_),
            .in1(N__5599),
            .in2(_gnd_net_),
            .in3(N__4726),
            .lcout(beamYZ0Z_8),
            .ltout(),
            .carryin(un21_beamy_cry_7),
            .carryout(un21_beamy_cry_8),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam beamY_9_LC_6_4_7.C_ON=1'b0;
    defparam beamY_9_LC_6_4_7.SEQ_MODE=4'b1000;
    defparam beamY_9_LC_6_4_7.LUT_INIT=16'b0001000100100010;
    LogicCell40 beamY_9_LC_6_4_7 (
            .in0(N__5628),
            .in1(N__5362),
            .in2(_gnd_net_),
            .in3(N__4816),
            .lcout(beamYZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7370),
            .ce(N__6250),
            .sr(_gnd_net_));
    defparam visibleY_2_LC_6_5_0.C_ON=1'b0;
    defparam visibleY_2_LC_6_5_0.SEQ_MODE=4'b1000;
    defparam visibleY_2_LC_6_5_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 visibleY_2_LC_6_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5535),
            .lcout(visibleYZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7365),
            .ce(N__7296),
            .sr(_gnd_net_));
    defparam TextOutputEnabled_LC_6_5_3.C_ON=1'b0;
    defparam TextOutputEnabled_LC_6_5_3.SEQ_MODE=4'b1000;
    defparam TextOutputEnabled_LC_6_5_3.LUT_INIT=16'b0100000000000000;
    LogicCell40 TextOutputEnabled_LC_6_5_3 (
            .in0(N__5161),
            .in1(N__4813),
            .in2(N__4804),
            .in3(N__4795),
            .lcout(TextOutputEnabledZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7365),
            .ce(N__7296),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_6_5.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_6_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_6_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_sbtinv_LC_6_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4942),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_7_0.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_7_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_7_0 (
            .in0(_gnd_net_),
            .in1(N__5807),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_7_0_),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSI_LC_6_7_1.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSI_LC_6_7_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSI_LC_6_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSI_LC_6_7_1 (
            .in0(_gnd_net_),
            .in1(N__4768),
            .in2(N__5028),
            .in3(N__4762),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2_c_RNILSVSIZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GT_LC_6_7_2.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GT_LC_6_7_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GT_LC_6_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GT_LC_6_7_2 (
            .in0(_gnd_net_),
            .in1(N__5022),
            .in2(N__4915),
            .in3(N__4759),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3_c_RNI3U4GTZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7C11_LC_6_7_3.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7C11_LC_6_7_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7C11_LC_6_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7C11_LC_6_7_3 (
            .in0(_gnd_net_),
            .in1(N__4897),
            .in2(N__5029),
            .in3(N__4756),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNI7H7CZ0Z11),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_6_7_4.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_6_7_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_6_7_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_inv_LC_6_7_4 (
            .in0(_gnd_net_),
            .in1(N__4858),
            .in2(N__4753),
            .in3(N__5023),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_i_7),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGC41_LC_6_7_5.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGC41_LC_6_7_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGC41_LC_6_7_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGC41_LC_6_7_5 (
            .in0(_gnd_net_),
            .in1(N__4834),
            .in2(_gnd_net_),
            .in3(N__4963),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41),
            .ltout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_cry_6_c_RNIRKGCZ0Z41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_3_LC_6_7_6.C_ON=1'b0;
    defparam Pixel_RNO_3_LC_6_7_6.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_3_LC_6_7_6.LUT_INIT=16'b1111101000001010;
    LogicCell40 Pixel_RNO_3_LC_6_7_6 (
            .in0(N__4957),
            .in1(_gnd_net_),
            .in2(N__4960),
            .in3(N__4948),
            .lcout(N_76),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_7_LC_6_7_7.C_ON=1'b0;
    defparam Pixel_RNO_7_LC_6_7_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_7_LC_6_7_7.LUT_INIT=16'b1111110100000010;
    LogicCell40 Pixel_RNO_7_LC_6_7_7 (
            .in0(N__5808),
            .in1(N__5842),
            .in2(N__5782),
            .in3(N__4956),
            .lcout(Pixel_RNOZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_8_0.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_8_0 (
            .in0(_gnd_net_),
            .in1(N__4941),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000B_LC_6_8_1.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000B_LC_6_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000B_LC_6_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000B_LC_6_8_1 (
            .in0(_gnd_net_),
            .in1(N__4883),
            .in2(N__4924),
            .in3(N__4906),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un61_sum_sbtinv_RNIP000BZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_2),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SE_LC_6_8_2.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SE_LC_6_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SE_LC_6_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SE_LC_6_8_2 (
            .in0(_gnd_net_),
            .in1(N__4903),
            .in2(N__4888),
            .in3(N__4891),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3_c_RNISH1SEZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_3),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OG_LC_6_8_3.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OG_LC_6_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OG_LC_6_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OG_LC_6_8_3 (
            .in0(_gnd_net_),
            .in1(N__4887),
            .in2(N__4867),
            .in3(N__4852),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNIS14OGZ0),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI2VO741_LC_6_8_4.C_ON=1'b1;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI2VO741_LC_6_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI2VO741_LC_6_8_4.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNI2VO741_LC_6_8_4 (
            .in0(N__5027),
            .in1(N__4849),
            .in2(N__4843),
            .in3(N__4828),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un75_sum_axb_7),
            .ltout(),
            .carryin(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBI_LC_6_8_5.C_ON=1'b0;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBI_LC_6_8_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBI_LC_6_8_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBI_LC_6_8_5 (
            .in0(_gnd_net_),
            .in1(N__4825),
            .in2(_gnd_net_),
            .in3(N__4819),
            .lcout(chessboardpixel_un32_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNIKDGBIZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIQCL_1_LC_6_8_7.C_ON=1'b0;
    defparam beamX_RNIQCL_1_LC_6_8_7.SEQ_MODE=4'b0000;
    defparam beamX_RNIQCL_1_LC_6_8_7.LUT_INIT=16'b0000011100001111;
    LogicCell40 beamX_RNIQCL_1_LC_6_8_7 (
            .in0(N__6344),
            .in1(N__6314),
            .in2(N__6649),
            .in3(N__6283),
            .lcout(un18_beamylt4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_0_c_LC_6_9_0.C_ON=1'b1;
    defparam un5_vx_cry_0_c_LC_6_9_0.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_0_c_LC_6_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un5_vx_cry_0_c_LC_6_9_0 (
            .in0(_gnd_net_),
            .in1(N__6281),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(un5_vx_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_1_LC_6_9_1.C_ON=1'b1;
    defparam beamX_1_LC_6_9_1.SEQ_MODE=4'b1000;
    defparam beamX_1_LC_6_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_1_LC_6_9_1 (
            .in0(N__6282),
            .in1(N__6313),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(beamXZ0Z_1),
            .ltout(),
            .carryin(un5_vx_cry_0),
            .carryout(un5_vx_cry_1),
            .clk(N__7358),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_1_c_RNIRP5_LC_6_9_2.C_ON=1'b1;
    defparam un5_vx_cry_1_c_RNIRP5_LC_6_9_2.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_1_c_RNIRP5_LC_6_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_vx_cry_1_c_RNIRP5_LC_6_9_2 (
            .in0(_gnd_net_),
            .in1(N__6343),
            .in2(_gnd_net_),
            .in3(N__5002),
            .lcout(c_if_generate_plus_mult1_un75_sum),
            .ltout(),
            .carryin(un5_vx_cry_1),
            .carryout(un5_vx_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_2_c_RNITS6_LC_6_9_3.C_ON=1'b1;
    defparam un5_vx_cry_2_c_RNITS6_LC_6_9_3.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_2_c_RNITS6_LC_6_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_vx_cry_2_c_RNITS6_LC_6_9_3 (
            .in0(_gnd_net_),
            .in1(N__6642),
            .in2(N__7782),
            .in3(N__4999),
            .lcout(c_if_generate_plus_mult1_un68_sum),
            .ltout(),
            .carryin(un5_vx_cry_2),
            .carryout(un5_vx_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_3_c_RNIVV7_LC_6_9_4.C_ON=1'b1;
    defparam un5_vx_cry_3_c_RNIVV7_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_3_c_RNIVV7_LC_6_9_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_vx_cry_3_c_RNIVV7_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(N__6710),
            .in2(_gnd_net_),
            .in3(N__4975),
            .lcout(c_if_generate_plus_mult1_un61_sum),
            .ltout(),
            .carryin(un5_vx_cry_3),
            .carryout(un5_vx_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_4_c_RNI139_LC_6_9_5.C_ON=1'b1;
    defparam un5_vx_cry_4_c_RNI139_LC_6_9_5.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_4_c_RNI139_LC_6_9_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_vx_cry_4_c_RNI139_LC_6_9_5 (
            .in0(_gnd_net_),
            .in1(N__6674),
            .in2(_gnd_net_),
            .in3(N__4972),
            .lcout(c_if_generate_plus_mult1_un47_sum1_0),
            .ltout(),
            .carryin(un5_vx_cry_4),
            .carryout(un5_vx_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_5_c_RNI36A_LC_6_9_6.C_ON=1'b1;
    defparam un5_vx_cry_5_c_RNI36A_LC_6_9_6.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_5_c_RNI36A_LC_6_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_vx_cry_5_c_RNI36A_LC_6_9_6 (
            .in0(_gnd_net_),
            .in1(N__7774),
            .in2(N__6748),
            .in3(N__4969),
            .lcout(c_if_generate_plus_mult1_un47_sum_1),
            .ltout(),
            .carryin(un5_vx_cry_5),
            .carryout(un5_vx_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_6_c_RNI59B_LC_6_9_7.C_ON=1'b1;
    defparam un5_vx_cry_6_c_RNI59B_LC_6_9_7.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_6_c_RNI59B_LC_6_9_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 un5_vx_cry_6_c_RNI59B_LC_6_9_7 (
            .in0(_gnd_net_),
            .in1(N__7135),
            .in2(_gnd_net_),
            .in3(N__4966),
            .lcout(un5_vx_cry_6_c_RNI59BZ0),
            .ltout(),
            .carryin(un5_vx_cry_6),
            .carryout(un5_vx_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_7_c_RNI7CC_LC_6_10_0.C_ON=1'b1;
    defparam un5_vx_cry_7_c_RNI7CC_LC_6_10_0.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_7_c_RNI7CC_LC_6_10_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 un5_vx_cry_7_c_RNI7CC_LC_6_10_0 (
            .in0(_gnd_net_),
            .in1(N__5899),
            .in2(N__7783),
            .in3(N__5062),
            .lcout(c_if_generate_plus_mult1_un47_sum_0_0),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(un5_vx_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_8_c_RNI9FD_LC_6_10_1.C_ON=1'b0;
    defparam un5_vx_cry_8_c_RNI9FD_LC_6_10_1.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_8_c_RNI9FD_LC_6_10_1.LUT_INIT=16'b1100110000110011;
    LogicCell40 un5_vx_cry_8_c_RNI9FD_LC_6_10_1 (
            .in0(_gnd_net_),
            .in1(N__5861),
            .in2(_gnd_net_),
            .in3(N__5059),
            .lcout(CO3_0),
            .ltout(CO3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TextOutputEnabled_RNO_3_LC_6_10_2.C_ON=1'b0;
    defparam TextOutputEnabled_RNO_3_LC_6_10_2.SEQ_MODE=4'b0000;
    defparam TextOutputEnabled_RNO_3_LC_6_10_2.LUT_INIT=16'b1100101000001010;
    LogicCell40 TextOutputEnabled_RNO_3_LC_6_10_2 (
            .in0(N__5988),
            .in1(N__6807),
            .in2(N__5056),
            .in3(N__6508),
            .lcout(N_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_7_c_RNIL451_LC_6_10_3.C_ON=1'b0;
    defparam un5_vx_cry_7_c_RNIL451_LC_6_10_3.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_7_c_RNIL451_LC_6_10_3.LUT_INIT=16'b0110011010011001;
    LogicCell40 un5_vx_cry_7_c_RNIL451_LC_6_10_3 (
            .in0(N__7439),
            .in1(N__6476),
            .in2(_gnd_net_),
            .in3(N__6027),
            .lcout(N_13_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_6_c_RNI59B_1_LC_6_10_4.C_ON=1'b0;
    defparam un5_vx_cry_6_c_RNI59B_1_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_6_c_RNI59B_1_LC_6_10_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 un5_vx_cry_6_c_RNI59B_1_LC_6_10_4 (
            .in0(N__6475),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(un5_vx_i_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_7_c_RNICLN_LC_6_10_5.C_ON=1'b0;
    defparam un5_vx_cry_7_c_RNICLN_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_7_c_RNICLN_LC_6_10_5.LUT_INIT=16'b0000000000110011;
    LogicCell40 un5_vx_cry_7_c_RNICLN_LC_6_10_5 (
            .in0(_gnd_net_),
            .in1(N__6474),
            .in2(_gnd_net_),
            .in3(N__6026),
            .lcout(N_3_0),
            .ltout(N_3_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_6_10_6.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_6_10_6.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_6_10_6.LUT_INIT=16'b0100011111001111;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx_LC_6_10_6 (
            .in0(N__6028),
            .in1(N__7440),
            .in2(N__5041),
            .in3(N__6479),
            .lcout(if_generate_plus_mult1_un47_sum_1_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_5_sbtinv_LC_6_10_7.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_5_sbtinv_LC_6_10_7.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_5_sbtinv_LC_6_10_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_axb_5_sbtinv_LC_6_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7435),
            .lcout(c_if_generate_plus_mult1_un47_sum_0_axb_5_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_11_0.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_11_0.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 c_if_generate_plus_mult1_un75_sum_cry_1_c_LC_6_11_0 (
            .in0(_gnd_net_),
            .in1(N__5038),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(c_if_generate_plus_mult1_un75_sum_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_11_1.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_11_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 c_if_generate_plus_mult1_un75_sum_cry_2_c_inv_LC_6_11_1 (
            .in0(_gnd_net_),
            .in1(N__5208),
            .in2(N__5128),
            .in3(N__5185),
            .lcout(G_253),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un75_sum_cry_1),
            .carryout(c_if_generate_plus_mult1_un75_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un75_sum_cry_3_c_LC_6_11_2.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un75_sum_cry_3_c_LC_6_11_2.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un75_sum_cry_3_c_LC_6_11_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 c_if_generate_plus_mult1_un75_sum_cry_3_c_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(N__5215),
            .in2(N__5191),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un75_sum_cry_2),
            .carryout(c_if_generate_plus_mult1_un75_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_11_3.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_11_3.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_11_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 c_if_generate_plus_mult1_un75_sum_cry_4_c_LC_6_11_3 (
            .in0(_gnd_net_),
            .in1(N__5209),
            .in2(N__5200),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un75_sum_cry_3),
            .carryout(c_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam TextOutputEnabled_RNO_1_LC_6_11_4.C_ON=1'b0;
    defparam TextOutputEnabled_RNO_1_LC_6_11_4.SEQ_MODE=4'b0000;
    defparam TextOutputEnabled_RNO_1_LC_6_11_4.LUT_INIT=16'b0000110100000111;
    LogicCell40 TextOutputEnabled_RNO_1_LC_6_11_4 (
            .in0(N__5189),
            .in1(N__5170),
            .in2(N__5119),
            .in3(N__5164),
            .lcout(un9_r_1lt6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un68_sum_i_LC_6_11_7.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un68_sum_i_LC_6_11_7.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un68_sum_i_LC_6_11_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 c_if_generate_plus_mult1_un68_sum_i_LC_6_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5150),
            .lcout(c_if_generate_plus_mult1_un68_sum_iZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un9_r_0lto3_sbtinv_LC_6_12_3.C_ON=1'b0;
    defparam un9_r_0lto3_sbtinv_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam un9_r_0lto3_sbtinv_LC_6_12_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un9_r_0lto3_sbtinv_LC_6_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5110),
            .lcout(un9_r_0lto3_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_N_404_i_LC_6_12_4.C_ON=1'b0;
    defparam c_N_404_i_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam c_N_404_i_LC_6_12_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 c_N_404_i_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5971),
            .lcout(N_404_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_6_12_7.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_6_12_7.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_6_12_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_sbtinv_5_LC_6_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6070),
            .lcout(c_if_generate_plus_mult1_un54_sum_i_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_0_LC_7_3_0.C_ON=1'b0;
    defparam beamY_0_LC_7_3_0.SEQ_MODE=4'b1000;
    defparam beamY_0_LC_7_3_0.LUT_INIT=16'b0001000110101010;
    LogicCell40 beamY_0_LC_7_3_0 (
            .in0(N__5336),
            .in1(N__5363),
            .in2(_gnd_net_),
            .in3(N__6249),
            .lcout(beamYZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7375),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_1_LC_7_3_3.C_ON=1'b0;
    defparam beamY_1_LC_7_3_3.SEQ_MODE=4'b1000;
    defparam beamY_1_LC_7_3_3.LUT_INIT=16'b0101001001110000;
    LogicCell40 beamY_1_LC_7_3_3 (
            .in0(N__6248),
            .in1(N__5364),
            .in2(N__5299),
            .in3(N__5337),
            .lcout(beamYZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7375),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI9DLC_2_LC_7_4_0.C_ON=1'b0;
    defparam beamY_RNI9DLC_2_LC_7_4_0.SEQ_MODE=4'b0000;
    defparam beamY_RNI9DLC_2_LC_7_4_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 beamY_RNI9DLC_2_LC_7_4_0 (
            .in0(N__5305),
            .in1(N__5533),
            .in2(N__5272),
            .in3(N__5314),
            .lcout(beamY_RNI9DLCZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIC725_0_LC_7_4_1.C_ON=1'b0;
    defparam beamY_RNIC725_0_LC_7_4_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIC725_0_LC_7_4_1.LUT_INIT=16'b0001000000000000;
    LogicCell40 beamY_RNIC725_0_LC_7_4_1 (
            .in0(N__5597),
            .in1(N__5335),
            .in2(N__5629),
            .in3(N__5444),
            .lcout(un5_beamx_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIN4H2_5_LC_7_4_2.C_ON=1'b0;
    defparam beamY_RNIN4H2_5_LC_7_4_2.SEQ_MODE=4'b0000;
    defparam beamY_RNIN4H2_5_LC_7_4_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNIN4H2_5_LC_7_4_2 (
            .in0(_gnd_net_),
            .in1(N__5678),
            .in2(_gnd_net_),
            .in3(N__5654),
            .lcout(un1_beamy_4),
            .ltout(un1_beamy_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIH3B6_7_LC_7_4_3.C_ON=1'b0;
    defparam beamY_RNIH3B6_7_LC_7_4_3.SEQ_MODE=4'b0000;
    defparam beamY_RNIH3B6_7_LC_7_4_3.LUT_INIT=16'b0000000011000000;
    LogicCell40 beamY_RNIH3B6_7_LC_7_4_3 (
            .in0(_gnd_net_),
            .in1(N__5256),
            .in2(N__5308),
            .in3(N__5565),
            .lcout(un8_beamylto9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNITAH2_9_LC_7_4_4.C_ON=1'b0;
    defparam beamY_RNITAH2_9_LC_7_4_4.SEQ_MODE=4'b0000;
    defparam beamY_RNITAH2_9_LC_7_4_4.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNITAH2_9_LC_7_4_4 (
            .in0(_gnd_net_),
            .in1(N__5623),
            .in2(_gnd_net_),
            .in3(N__5596),
            .lcout(un8_beamy_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIEIP3_1_LC_7_4_5.C_ON=1'b0;
    defparam beamY_RNIEIP3_1_LC_7_4_5.SEQ_MODE=4'b0000;
    defparam beamY_RNIEIP3_1_LC_7_4_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 beamY_RNIEIP3_1_LC_7_4_5 (
            .in0(N__5489),
            .in1(N__5566),
            .in2(_gnd_net_),
            .in3(N__5294),
            .lcout(un5_beamx_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_RNO_0_LC_7_4_6.C_ON=1'b0;
    defparam VSync_1_RNO_0_LC_7_4_6.SEQ_MODE=4'b0000;
    defparam VSync_1_RNO_0_LC_7_4_6.LUT_INIT=16'b0000000100000011;
    LogicCell40 VSync_1_RNO_0_LC_7_4_6 (
            .in0(N__5295),
            .in1(N__5569),
            .in2(N__5449),
            .in3(N__5534),
            .lcout(),
            .ltout(un1_beamylto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam VSync_1_LC_7_4_7.C_ON=1'b0;
    defparam VSync_1_LC_7_4_7.SEQ_MODE=4'b1000;
    defparam VSync_1_LC_7_4_7.LUT_INIT=16'b1111111101111111;
    LogicCell40 VSync_1_LC_7_4_7 (
            .in0(N__5271),
            .in1(N__5257),
            .in2(N__5248),
            .in3(N__5491),
            .lcout(VSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7373),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNIHUG2_3_LC_7_5_1.C_ON=1'b0;
    defparam beamY_RNIHUG2_3_LC_7_5_1.SEQ_MODE=4'b0000;
    defparam beamY_RNIHUG2_3_LC_7_5_1.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamY_RNIHUG2_3_LC_7_5_1 (
            .in0(_gnd_net_),
            .in1(N__5442),
            .in2(_gnd_net_),
            .in3(N__5527),
            .lcout(),
            .ltout(un4_beamylt6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNI2KA6_5_LC_7_5_2.C_ON=1'b0;
    defparam beamY_RNI2KA6_5_LC_7_5_2.SEQ_MODE=4'b0000;
    defparam beamY_RNI2KA6_5_LC_7_5_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 beamY_RNI2KA6_5_LC_7_5_2 (
            .in0(N__5679),
            .in1(N__5655),
            .in2(N__5632),
            .in3(N__5487),
            .lcout(),
            .ltout(un4_beamylt8_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_9_LC_7_5_3.C_ON=1'b0;
    defparam beamY_RNISI4A_9_LC_7_5_3.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_9_LC_7_5_3.LUT_INIT=16'b1010101010101000;
    LogicCell40 beamY_RNISI4A_9_LC_7_5_3 (
            .in0(N__5627),
            .in1(N__5598),
            .in2(N__5572),
            .in3(N__5567),
            .lcout(un4_beamy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamY_RNISI4A_3_LC_7_5_6.C_ON=1'b0;
    defparam beamY_RNISI4A_3_LC_7_5_6.SEQ_MODE=4'b0000;
    defparam beamY_RNISI4A_3_LC_7_5_6.LUT_INIT=16'b0111000011110000;
    LogicCell40 beamY_RNISI4A_3_LC_7_5_6 (
            .in0(N__5528),
            .in1(N__5488),
            .in2(N__5458),
            .in3(N__5443),
            .lcout(un8_beamy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_5_LC_7_6_0.C_ON=1'b0;
    defparam Pixel_RNO_5_LC_7_6_0.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_5_LC_7_6_0.LUT_INIT=16'b1011111111111111;
    LogicCell40 Pixel_RNO_5_LC_7_6_0 (
            .in0(N__5806),
            .in1(N__5840),
            .in2(N__5827),
            .in3(N__5781),
            .lcout(),
            .ltout(Pixel_RNOZ0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_1_LC_7_6_1.C_ON=1'b0;
    defparam Pixel_RNO_1_LC_7_6_1.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_1_LC_7_6_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 Pixel_RNO_1_LC_7_6_1 (
            .in0(_gnd_net_),
            .in1(N__5413),
            .in2(N__5407),
            .in3(N__5761),
            .lcout(),
            .ltout(N_45_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_0_LC_7_6_2.C_ON=1'b0;
    defparam Pixel_RNO_0_LC_7_6_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_0_LC_7_6_2.LUT_INIT=16'b0100010010110100;
    LogicCell40 Pixel_RNO_0_LC_7_6_2 (
            .in0(N__6361),
            .in1(N__6415),
            .in2(N__5404),
            .in3(N__5401),
            .lcout(),
            .ltout(N_74_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PixelZ0_LC_7_6_3.C_ON=1'b0;
    defparam PixelZ0_LC_7_6_3.SEQ_MODE=4'b1000;
    defparam PixelZ0_LC_7_6_3.LUT_INIT=16'b1011100000000000;
    LogicCell40 PixelZ0_LC_7_6_3 (
            .in0(N__7546),
            .in1(N__5395),
            .in2(N__5389),
            .in3(N__5752),
            .lcout(Pixel_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVPixelZ0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_6_LC_7_6_7.C_ON=1'b0;
    defparam Pixel_RNO_6_LC_7_6_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_6_LC_7_6_7.LUT_INIT=16'b1111111110111111;
    LogicCell40 Pixel_RNO_6_LC_7_6_7 (
            .in0(N__5841),
            .in1(N__5823),
            .in2(N__5809),
            .in3(N__5780),
            .lcout(Pixel_RNOZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI8P51_4_LC_7_7_0.C_ON=1'b0;
    defparam beamX_RNI8P51_4_LC_7_7_0.SEQ_MODE=4'b0000;
    defparam beamX_RNI8P51_4_LC_7_7_0.LUT_INIT=16'b0011001100010011;
    LogicCell40 beamX_RNI8P51_4_LC_7_7_0 (
            .in0(N__6712),
            .in1(N__6743),
            .in2(N__6684),
            .in3(N__5746),
            .lcout(un13_beamylt7),
            .ltout(un13_beamylt7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutputEnabled_LC_7_7_1.C_ON=1'b0;
    defparam OutputEnabled_LC_7_7_1.SEQ_MODE=4'b1000;
    defparam OutputEnabled_LC_7_7_1.LUT_INIT=16'b0011101100000000;
    LogicCell40 OutputEnabled_LC_7_7_1 (
            .in0(N__7138),
            .in1(N__7166),
            .in2(N__5755),
            .in3(N__5710),
            .lcout(OutputEnabledZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7360),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIR4B_9_LC_7_7_3.C_ON=1'b0;
    defparam beamX_RNIR4B_9_LC_7_7_3.SEQ_MODE=4'b0000;
    defparam beamX_RNIR4B_9_LC_7_7_3.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_RNIR4B_9_LC_7_7_3 (
            .in0(_gnd_net_),
            .in1(N__5871),
            .in2(_gnd_net_),
            .in3(N__5897),
            .lcout(un1_beamx_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNII5M_9_LC_7_7_4.C_ON=1'b0;
    defparam beamX_RNII5M_9_LC_7_7_4.SEQ_MODE=4'b0000;
    defparam beamX_RNII5M_9_LC_7_7_4.LUT_INIT=16'b1000000000000000;
    LogicCell40 beamX_RNII5M_9_LC_7_7_4 (
            .in0(N__5896),
            .in1(N__7136),
            .in2(N__5872),
            .in3(N__6744),
            .lcout(),
            .ltout(un18_beamylto9_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIVEM1_4_LC_7_7_5.C_ON=1'b0;
    defparam beamX_RNIVEM1_4_LC_7_7_5.SEQ_MODE=4'b0000;
    defparam beamX_RNIVEM1_4_LC_7_7_5.LUT_INIT=16'b1101000011000000;
    LogicCell40 beamX_RNIVEM1_4_LC_7_7_5 (
            .in0(N__5745),
            .in1(N__6678),
            .in2(N__5734),
            .in3(N__6711),
            .lcout(),
            .ltout(un18_beamylt10_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIT9ER_10_LC_7_7_6.C_ON=1'b0;
    defparam beamX_RNIT9ER_10_LC_7_7_6.SEQ_MODE=4'b0000;
    defparam beamX_RNIT9ER_10_LC_7_7_6.LUT_INIT=16'b0000000000000001;
    LogicCell40 beamX_RNIT9ER_10_LC_7_7_6 (
            .in0(N__5731),
            .in1(N__7205),
            .in2(N__5722),
            .in3(N__5719),
            .lcout(un15_beamy_2),
            .ltout(un15_beamy_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNISO4T_7_LC_7_7_7.C_ON=1'b0;
    defparam beamX_RNISO4T_7_LC_7_7_7.SEQ_MODE=4'b0000;
    defparam beamX_RNISO4T_7_LC_7_7_7.LUT_INIT=16'b0010000011110000;
    LogicCell40 beamX_RNISO4T_7_LC_7_7_7 (
            .in0(N__7137),
            .in1(N__5704),
            .in2(N__5698),
            .in3(N__7165),
            .lcout(beamX_RNISO4TZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un8_beamx_cry_1_c_LC_7_8_0.C_ON=1'b1;
    defparam un8_beamx_cry_1_c_LC_7_8_0.SEQ_MODE=4'b0000;
    defparam un8_beamx_cry_1_c_LC_7_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 un8_beamx_cry_1_c_LC_7_8_0 (
            .in0(_gnd_net_),
            .in1(N__6318),
            .in2(N__6289),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(un8_beamx_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_2_LC_7_8_1.C_ON=1'b1;
    defparam beamX_2_LC_7_8_1.SEQ_MODE=4'b1000;
    defparam beamX_2_LC_7_8_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_2_LC_7_8_1 (
            .in0(_gnd_net_),
            .in1(N__6346),
            .in2(_gnd_net_),
            .in3(N__5917),
            .lcout(beamXZ0Z_2),
            .ltout(),
            .carryin(un8_beamx_cry_1),
            .carryout(un8_beamx_cry_2),
            .clk(N__7355),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_3_LC_7_8_2.C_ON=1'b1;
    defparam beamX_3_LC_7_8_2.SEQ_MODE=4'b1000;
    defparam beamX_3_LC_7_8_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_3_LC_7_8_2 (
            .in0(_gnd_net_),
            .in1(N__6648),
            .in2(_gnd_net_),
            .in3(N__5914),
            .lcout(beamXZ0Z_3),
            .ltout(),
            .carryin(un8_beamx_cry_2),
            .carryout(un8_beamx_cry_3),
            .clk(N__7355),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_4_LC_7_8_3.C_ON=1'b1;
    defparam beamX_4_LC_7_8_3.SEQ_MODE=4'b1000;
    defparam beamX_4_LC_7_8_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_4_LC_7_8_3 (
            .in0(N__6239),
            .in1(N__6715),
            .in2(_gnd_net_),
            .in3(N__5911),
            .lcout(beamXZ0Z_4),
            .ltout(),
            .carryin(un8_beamx_cry_3),
            .carryout(un8_beamx_cry_4),
            .clk(N__7355),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_5_LC_7_8_4.C_ON=1'b1;
    defparam beamX_5_LC_7_8_4.SEQ_MODE=4'b1000;
    defparam beamX_5_LC_7_8_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_5_LC_7_8_4 (
            .in0(_gnd_net_),
            .in1(N__6683),
            .in2(_gnd_net_),
            .in3(N__5908),
            .lcout(beamXZ0Z_5),
            .ltout(),
            .carryin(un8_beamx_cry_4),
            .carryout(un8_beamx_cry_5),
            .clk(N__7355),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_6_LC_7_8_5.C_ON=1'b1;
    defparam beamX_6_LC_7_8_5.SEQ_MODE=4'b1000;
    defparam beamX_6_LC_7_8_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_6_LC_7_8_5 (
            .in0(_gnd_net_),
            .in1(N__6747),
            .in2(_gnd_net_),
            .in3(N__5905),
            .lcout(beamXZ0Z_6),
            .ltout(),
            .carryin(un8_beamx_cry_5),
            .carryout(un8_beamx_cry_6),
            .clk(N__7355),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_7_LC_7_8_6.C_ON=1'b1;
    defparam beamX_7_LC_7_8_6.SEQ_MODE=4'b1000;
    defparam beamX_7_LC_7_8_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_7_LC_7_8_6 (
            .in0(_gnd_net_),
            .in1(N__7140),
            .in2(_gnd_net_),
            .in3(N__5902),
            .lcout(beamXZ0Z_7),
            .ltout(),
            .carryin(un8_beamx_cry_6),
            .carryout(un8_beamx_cry_7),
            .clk(N__7355),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_8_LC_7_8_7.C_ON=1'b1;
    defparam beamX_8_LC_7_8_7.SEQ_MODE=4'b1000;
    defparam beamX_8_LC_7_8_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_8_LC_7_8_7 (
            .in0(_gnd_net_),
            .in1(N__5898),
            .in2(_gnd_net_),
            .in3(N__5875),
            .lcout(beamXZ0Z_8),
            .ltout(),
            .carryin(un8_beamx_cry_7),
            .carryout(un8_beamx_cry_8),
            .clk(N__7355),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_9_LC_7_9_0.C_ON=1'b1;
    defparam beamX_9_LC_7_9_0.SEQ_MODE=4'b1000;
    defparam beamX_9_LC_7_9_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 beamX_9_LC_7_9_0 (
            .in0(_gnd_net_),
            .in1(N__5867),
            .in2(_gnd_net_),
            .in3(N__5845),
            .lcout(beamXZ0Z_9),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(un8_beamx_cry_9),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_10_LC_7_9_1.C_ON=1'b0;
    defparam beamX_10_LC_7_9_1.SEQ_MODE=4'b1000;
    defparam beamX_10_LC_7_9_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 beamX_10_LC_7_9_1 (
            .in0(N__6234),
            .in1(N__7204),
            .in2(_gnd_net_),
            .in3(N__5953),
            .lcout(beamXZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_0_LC_7_9_2.C_ON=1'b0;
    defparam beamX_0_LC_7_9_2.SEQ_MODE=4'b1000;
    defparam beamX_0_LC_7_9_2.LUT_INIT=16'b0000000000110011;
    LogicCell40 beamX_0_LC_7_9_2 (
            .in0(_gnd_net_),
            .in1(N__6235),
            .in2(_gnd_net_),
            .in3(N__6288),
            .lcout(un5_vx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7361),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_6_c_RNI59B_0_LC_7_9_3.C_ON=1'b0;
    defparam un5_vx_cry_6_c_RNI59B_0_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_6_c_RNI59B_0_LC_7_9_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 un5_vx_cry_6_c_RNI59B_0_LC_7_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6477),
            .lcout(un5_vx_i_25),
            .ltout(un5_vx_i_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_7_9_4.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_7_9_4.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_7_9_4.LUT_INIT=16'b0000111111110000;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx_LC_7_9_4 (
            .in0(N__7438),
            .in1(N__6803),
            .in2(N__5950),
            .in3(N__6029),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_3_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_9_5.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_9_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_cry_3_ma_LC_7_9_5 (
            .in0(N__6801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7436),
            .lcout(if_generate_plus_mult1_un47_sum_0_cry_3_ma),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_9_6.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_9_6.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_9_6.LUT_INIT=16'b0011001111111111;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx_LC_7_9_6 (
            .in0(N__6478),
            .in1(N__7434),
            .in2(_gnd_net_),
            .in3(N__6800),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_2_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un5_vx_cry_8_c_RNIL451_LC_7_9_7.C_ON=1'b0;
    defparam un5_vx_cry_8_c_RNIL451_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_8_c_RNIL451_LC_7_9_7.LUT_INIT=16'b0101010111111111;
    LogicCell40 un5_vx_cry_8_c_RNIL451_LC_7_9_7 (
            .in0(N__6802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7437),
            .lcout(N_186_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_10_0.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_1_cry_1_c_LC_7_10_0 (
            .in0(_gnd_net_),
            .in1(N__6610),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(c_if_generate_plus_mult1_un47_sum_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_m_2_LC_7_10_1.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un47_sum_m_2_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_m_2_LC_7_10_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_m_2_LC_7_10_1 (
            .in0(N__6574),
            .in1(N__7449),
            .in2(N__5947),
            .in3(N__5938),
            .lcout(if_generate_plus_mult1_un47_sum_m_2),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un47_sum_1_cry_1),
            .carryout(c_if_generate_plus_mult1_un47_sum_1_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_10_2.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_1_cry_3_s_LC_7_10_2 (
            .in0(_gnd_net_),
            .in1(N__5935),
            .in2(N__5929),
            .in3(N__5920),
            .lcout(c_if_generate_plus_mult1_un47_sum1_3),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un47_sum_1_cry_2),
            .carryout(c_if_generate_plus_mult1_un47_sum_1_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_10_3.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_1_cry_4_s_LC_7_10_3 (
            .in0(_gnd_net_),
            .in1(N__6046),
            .in2(N__7466),
            .in3(N__6040),
            .lcout(c_if_generate_plus_mult1_un47_sum1_4),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un47_sum_1_cry_3),
            .carryout(c_if_generate_plus_mult1_un47_sum_1_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_10_4.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_10_4.LUT_INIT=16'b1000000001111111;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_1_s_5_LC_7_10_4 (
            .in0(N__7450),
            .in1(N__6480),
            .in2(N__6034),
            .in3(N__6037),
            .lcout(c_if_generate_plus_mult1_un47_sum1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_8_LC_7_10_6.C_ON=1'b0;
    defparam visibleX_8_LC_7_10_6.SEQ_MODE=4'b1000;
    defparam visibleX_8_LC_7_10_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 visibleX_8_LC_7_10_6 (
            .in0(N__6033),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(visibleXZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7366),
            .ce(N__7294),
            .sr(_gnd_net_));
    defparam un5_vx_cry_8_c_RNI24IE_LC_7_11_0.C_ON=1'b0;
    defparam un5_vx_cry_8_c_RNI24IE_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam un5_vx_cry_8_c_RNI24IE_LC_7_11_0.LUT_INIT=16'b0001000110111011;
    LogicCell40 un5_vx_cry_8_c_RNI24IE_LC_7_11_0 (
            .in0(N__7454),
            .in1(N__5984),
            .in2(_gnd_net_),
            .in3(N__6503),
            .lcout(N_18),
            .ltout(N_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_axb_5_LC_7_11_1.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un54_sum_axb_5_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_axb_5_LC_7_11_1.LUT_INIT=16'b0011110001011010;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_axb_5_LC_7_11_1 (
            .in0(N__6004),
            .in1(N__6523),
            .in2(N__5998),
            .in3(N__7458),
            .lcout(c_if_generate_plus_mult1_un54_sum_axbZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_7_11_2.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_7_11_2.LUT_INIT=16'b0010001001110111;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_axb_2_l_fx_LC_7_11_2 (
            .in0(N__7455),
            .in1(N__6618),
            .in2(N__6141),
            .in3(N__6619),
            .lcout(if_generate_plus_mult1_un54_sum_axb_2_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_11_3.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_11_3.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_11_3.LUT_INIT=16'b1110111000100010;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_axb_4_l_fx_LC_7_11_3 (
            .in0(N__5995),
            .in1(N__7457),
            .in2(N__6142),
            .in3(N__6544),
            .lcout(if_generate_plus_mult1_un54_sum_axb_4_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_7_11_7.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_7_11_7.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_7_11_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_axb_3_l_fx_LC_7_11_7 (
            .in0(N__6504),
            .in1(N__6171),
            .in2(N__5989),
            .in3(N__7456),
            .lcout(if_generate_plus_mult1_un54_sum_axb_3_l_fx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_5_LC_7_12_0.C_ON=1'b1;
    defparam visibleX_5_LC_7_12_0.SEQ_MODE=4'b1000;
    defparam visibleX_5_LC_7_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleX_5_LC_7_12_0 (
            .in0(_gnd_net_),
            .in1(N__5969),
            .in2(_gnd_net_),
            .in3(N__5970),
            .lcout(visibleXZ0Z_5),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(c_if_generate_plus_mult1_un54_sum_cry_1),
            .clk(N__7372),
            .ce(N__7297),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_cry_2_s_LC_7_12_1 (
            .in0(_gnd_net_),
            .in1(N__6133),
            .in2(N__6205),
            .in3(N__6184),
            .lcout(if_generate_plus_mult1_un54_sum_cry_2_s),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un54_sum_cry_1),
            .carryout(c_if_generate_plus_mult1_un54_sum_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_12_2 (
            .in0(_gnd_net_),
            .in1(N__6181),
            .in2(N__6175),
            .in3(N__6145),
            .lcout(if_generate_plus_mult1_un54_sum_cry_3_s),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un54_sum_cry_2),
            .carryout(c_if_generate_plus_mult1_un54_sum_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 c_if_generate_plus_mult1_un61_sum_axb_5_LC_7_12_3 (
            .in0(N__6071),
            .in1(N__6134),
            .in2(N__6115),
            .in3(N__6097),
            .lcout(c_if_generate_plus_mult1_un61_sum_axbZ0Z_5),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un54_sum_cry_3),
            .carryout(c_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 c_if_generate_plus_mult1_un54_sum_s_5_LC_7_12_4 (
            .in0(_gnd_net_),
            .in1(N__6094),
            .in2(_gnd_net_),
            .in3(N__6088),
            .lcout(if_generate_plus_mult1_un54_sum_s_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_8_4_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_4_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_4_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_4_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_8_7_0.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_8_7_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_8_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_LC_8_7_0 (
            .in0(_gnd_net_),
            .in1(N__6386),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HC_LC_8_7_1.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HC_LC_8_7_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HC_LC_8_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HC_LC_8_7_1 (
            .in0(_gnd_net_),
            .in1(N__6441),
            .in2(N__6355),
            .in3(N__6052),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4_c_RNIQ0HCZ0),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_4),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_8_LC_8_7_2.C_ON=1'b1;
    defparam Pixel_RNO_8_LC_8_7_2.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_8_LC_8_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 Pixel_RNO_8_LC_8_7_2 (
            .in0(_gnd_net_),
            .in1(N__6886),
            .in2(N__6850),
            .in3(N__6049),
            .lcout(Pixel_RNOZ0Z_8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_5),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_8_7_3.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_8_7_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_8_7_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_inv_LC_8_7_3 (
            .in0(_gnd_net_),
            .in1(N__6442),
            .in2(N__6874),
            .in3(N__6845),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i_8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_6),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53L_LC_8_7_4.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53L_LC_8_7_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53L_LC_8_7_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53L_LC_8_7_4 (
            .in0(_gnd_net_),
            .in1(N__6862),
            .in2(_gnd_net_),
            .in3(N__6433),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0),
            .ltout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_cry_7_c_RNICN53LZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_2_LC_8_7_5.C_ON=1'b0;
    defparam Pixel_RNO_2_LC_8_7_5.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_2_LC_8_7_5.LUT_INIT=16'b0101001010111111;
    LogicCell40 Pixel_RNO_2_LC_8_7_5 (
            .in0(N__6387),
            .in1(N__6430),
            .in2(N__6418),
            .in3(N__6408),
            .lcout(N_53),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam Pixel_RNO_4_LC_8_7_7.C_ON=1'b0;
    defparam Pixel_RNO_4_LC_8_7_7.SEQ_MODE=4'b0000;
    defparam Pixel_RNO_4_LC_8_7_7.LUT_INIT=16'b0011100111001100;
    LogicCell40 Pixel_RNO_4_LC_8_7_7 (
            .in0(N__6409),
            .in1(N__6397),
            .in2(N__6391),
            .in3(N__6367),
            .lcout(N_81),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_RNIJK0C_5_LC_8_8_1.C_ON=1'b0;
    defparam visibleX_RNIJK0C_5_LC_8_8_1.SEQ_MODE=4'b0000;
    defparam visibleX_RNIJK0C_5_LC_8_8_1.LUT_INIT=16'b0011001100110011;
    LogicCell40 visibleX_RNIJK0C_5_LC_8_8_1 (
            .in0(_gnd_net_),
            .in1(N__6904),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNICPU5_10_LC_8_8_2.C_ON=1'b0;
    defparam beamX_RNICPU5_10_LC_8_8_2.SEQ_MODE=4'b0000;
    defparam beamX_RNICPU5_10_LC_8_8_2.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNICPU5_10_LC_8_8_2 (
            .in0(N__6713),
            .in1(N__6345),
            .in2(N__7206),
            .in3(N__6322),
            .lcout(),
            .ltout(un3_beamx_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNIKVE6_0_LC_8_8_3.C_ON=1'b0;
    defparam beamX_RNIKVE6_0_LC_8_8_3.SEQ_MODE=4'b0000;
    defparam beamX_RNIKVE6_0_LC_8_8_3.LUT_INIT=16'b0000000000010000;
    LogicCell40 beamX_RNIKVE6_0_LC_8_8_3 (
            .in0(N__6745),
            .in1(N__6646),
            .in2(N__6292),
            .in3(N__6284),
            .lcout(),
            .ltout(un3_beamx_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam beamX_RNI5457_5_LC_8_8_4.C_ON=1'b0;
    defparam beamX_RNI5457_5_LC_8_8_4.SEQ_MODE=4'b0000;
    defparam beamX_RNI5457_5_LC_8_8_4.LUT_INIT=16'b0000000000100000;
    LogicCell40 beamX_RNI5457_5_LC_8_8_4 (
            .in0(N__7167),
            .in1(N__7139),
            .in2(N__6253),
            .in3(N__6679),
            .lcout(beamX_RNI5457Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_RNO_0_LC_8_8_7.C_ON=1'b0;
    defparam HSync_1_RNO_0_LC_8_8_7.SEQ_MODE=4'b0000;
    defparam HSync_1_RNO_0_LC_8_8_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 HSync_1_RNO_0_LC_8_8_7 (
            .in0(N__6746),
            .in1(N__6714),
            .in2(N__6685),
            .in3(N__6647),
            .lcout(un1_beamxlt10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_6_LC_8_9_0.C_ON=1'b1;
    defparam visibleX_6_LC_8_9_0.SEQ_MODE=4'b1000;
    defparam visibleX_6_LC_8_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleX_6_LC_8_9_0 (
            .in0(_gnd_net_),
            .in1(N__6616),
            .in2(_gnd_net_),
            .in3(N__6617),
            .lcout(visibleXZ0Z_6),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(c_if_generate_plus_mult1_un47_sum_0_cry_1),
            .clk(N__7368),
            .ce(N__7291),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_9_1.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_9_1.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_cry_2_s_LC_8_9_1 (
            .in0(_gnd_net_),
            .in1(N__6589),
            .in2(N__6583),
            .in3(N__6562),
            .lcout(c_if_generate_plus_mult1_un47_sum0_2),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un47_sum_0_cry_1),
            .carryout(c_if_generate_plus_mult1_un47_sum_0_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_9_2.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_9_2.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_cry_3_0_s_LC_8_9_2 (
            .in0(_gnd_net_),
            .in1(N__6559),
            .in2(N__6553),
            .in3(N__6535),
            .lcout(c_if_generate_plus_mult1_un47_sum0_3),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un47_sum_0_cry_2),
            .carryout(c_if_generate_plus_mult1_un47_sum_0_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_9_3.C_ON=1'b1;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_9_3.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_cry_4_s_LC_8_9_3 (
            .in0(_gnd_net_),
            .in1(N__6778),
            .in2(N__6532),
            .in3(N__6514),
            .lcout(c_if_generate_plus_mult1_un47_sum0_4),
            .ltout(),
            .carryin(c_if_generate_plus_mult1_un47_sum_0_cry_3),
            .carryout(c_if_generate_plus_mult1_un47_sum_0_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_9_4.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_s_5_LC_8_9_4 (
            .in0(_gnd_net_),
            .in1(N__7467),
            .in2(_gnd_net_),
            .in3(N__6511),
            .lcout(c_if_generate_plus_mult1_un47_sum0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_7_LC_8_9_7.C_ON=1'b0;
    defparam visibleX_7_LC_8_9_7.SEQ_MODE=4'b1000;
    defparam visibleX_7_LC_8_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleX_7_LC_8_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6484),
            .lcout(visibleXZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7368),
            .ce(N__7291),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_10_0.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_LC_8_10_0 (
            .in0(_gnd_net_),
            .in1(N__7488),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BD1_LC_8_10_1.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BD1_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BD1_LC_8_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BD1_LC_8_10_1 (
            .in0(_gnd_net_),
            .in1(N__6912),
            .in2(N__6817),
            .in3(N__6832),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4_c_RNI91BDZ0Z1),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_4),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMK642_LC_8_10_2.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMK642_LC_8_10_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMK642_LC_8_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMK642_LC_8_10_2 (
            .in0(_gnd_net_),
            .in1(N__6928),
            .in2(N__6760),
            .in3(N__6829),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5_c_RNIMKZ0Z642),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_5),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3O524_LC_8_10_3.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3O524_LC_8_10_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3O524_LC_8_10_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6_c_RNI3O524_LC_8_10_3 (
            .in0(N__7041),
            .in1(N__6913),
            .in2(N__6952),
            .in3(N__6826),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_6),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_LC_8_10_4.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_LC_8_10_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_LC_8_10_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_LC_8_10_4 (
            .in0(_gnd_net_),
            .in1(N__6940),
            .in2(_gnd_net_),
            .in3(N__6823),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412),
            .ltout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3FZ0Z412_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_0_LC_8_10_5.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_0_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_0_LC_8_10_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_cry_7_c_RNI3F412_0_LC_8_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6820),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_RNIMN0C_8_LC_8_10_6.C_ON=1'b0;
    defparam visibleX_RNIMN0C_8_LC_8_10_6.SEQ_MODE=4'b0000;
    defparam visibleX_RNIMN0C_8_LC_8_10_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 visibleX_RNIMN0C_8_LC_8_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6772),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_10_7.C_ON=1'b0;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam c_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_10_7.LUT_INIT=16'b1010101001010101;
    LogicCell40 c_if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx_LC_8_10_7 (
            .in0(N__7459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6808),
            .lcout(if_generate_plus_mult1_un47_sum_0_axb_4_l_ofx),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_11_0.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_LC_8_11_0 (
            .in0(_gnd_net_),
            .in1(N__6771),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29R21_LC_8_11_1.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29R21_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29R21_LC_8_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29R21_LC_8_11_1 (
            .in0(_gnd_net_),
            .in1(N__7566),
            .in2(N__7792),
            .in3(N__6751),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4_c_RNI29RZ0Z21),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_4),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKV_LC_8_11_2.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKV_LC_8_11_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKV_LC_8_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKV_LC_8_11_2 (
            .in0(_gnd_net_),
            .in1(N__7578),
            .in2(N__7252),
            .in3(N__6943),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5_c_RNIBRKVZ0),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_5),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIS2GV1_LC_8_11_3.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIS2GV1_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIS2GV1_LC_8_11_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6_c_RNIS2GV1_LC_8_11_3 (
            .in0(N__6927),
            .in1(N__7567),
            .in2(N__7240),
            .in3(N__6934),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_6),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_LC_8_11_4.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_LC_8_11_4.LUT_INIT=16'b0110011010011001;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_LC_8_11_4 (
            .in0(N__7228),
            .in1(N__7579),
            .in2(_gnd_net_),
            .in3(N__6931),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PVZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_0_LC_8_11_6.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_0_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_0_LC_8_11_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_cry_7_c_RNIF3PV_0_LC_8_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6926),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un47_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_8_0.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_8_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_LC_9_8_0 (
            .in0(_gnd_net_),
            .in1(N__6903),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56B05_LC_9_8_1.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56B05_LC_9_8_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56B05_LC_9_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56B05_LC_9_8_1 (
            .in0(_gnd_net_),
            .in1(N__7495),
            .in2(N__7072),
            .in3(N__6877),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4_c_RNI56BZ0Z05),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_4),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIC7997_LC_9_8_2.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIC7997_LC_9_8_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIC7997_LC_9_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNIC7997_LC_9_8_2 (
            .in0(_gnd_net_),
            .in1(N__7051),
            .in2(N__6970),
            .in3(N__6865),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5_c_RNICZ0Z7997),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_5),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI25I2L_LC_9_8_3.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI25I2L_LC_9_8_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI25I2L_LC_9_8_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6_c_RNI25I2L_LC_9_8_3 (
            .in0(N__6849),
            .in1(N__7216),
            .in2(N__7021),
            .in3(N__6856),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un75_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_6),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJ19_LC_9_8_4.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJ19_LC_9_8_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJ19_LC_9_8_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJ19_LC_9_8_4 (
            .in0(_gnd_net_),
            .in1(N__6988),
            .in2(_gnd_net_),
            .in3(N__6853),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_cry_7_c_RNIHDJZ0Z19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEA08_LC_9_8_5.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEA08_LC_9_8_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEA08_LC_9_8_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEA08_LC_9_8_5 (
            .in0(N__7020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6965),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNINEAZ0Z08),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam HSync_1_LC_9_8_6.C_ON=1'b0;
    defparam HSync_1_LC_9_8_6.SEQ_MODE=4'b1000;
    defparam HSync_1_LC_9_8_6.LUT_INIT=16'b1111111111111011;
    LogicCell40 HSync_1_LC_9_8_6 (
            .in0(N__7210),
            .in1(N__7174),
            .in2(N__7147),
            .in3(N__7105),
            .lcout(HSync_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7362),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_RNIKL0C_6_LC_9_8_7.C_ON=1'b0;
    defparam visibleX_RNIKL0C_6_LC_9_8_7.SEQ_MODE=4'b0000;
    defparam visibleX_RNIKL0C_6_LC_9_8_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 visibleX_RNIKL0C_6_LC_9_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7063),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_9_0.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_9_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_LC_9_9_0 (
            .in0(_gnd_net_),
            .in1(N__7062),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTK2_LC_9_9_1.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTK2_LC_9_9_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTK2_LC_9_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTK2_LC_9_9_1 (
            .in0(_gnd_net_),
            .in1(N__7005),
            .in2(N__7477),
            .in3(N__7045),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4_c_RNIQKTKZ0Z2),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_4),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19M3_LC_9_9_2.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19M3_LC_9_9_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19M3_LC_9_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19M3_LC_9_9_2 (
            .in0(_gnd_net_),
            .in1(N__7042),
            .in2(N__7030),
            .in3(N__7009),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5_c_RNIF19MZ0Z3),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_5),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNI547N8_LC_9_9_3.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNI547N8_LC_9_9_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNI547N8_LC_9_9_3.LUT_INIT=16'b1001011001101001;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6_c_RNI547N8_LC_9_9_3 (
            .in0(N__6969),
            .in1(N__7006),
            .in2(N__6997),
            .in3(N__6982),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un68_sum_axb_8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_6),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_LC_9_9_4.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_LC_9_9_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_LC_9_9_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_LC_9_9_4 (
            .in0(_gnd_net_),
            .in1(N__6979),
            .in2(_gnd_net_),
            .in3(N__6973),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4),
            .ltout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1AZ0Z4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_0_LC_9_9_5.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_0_LC_9_9_5.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_0_LC_9_9_5.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_cry_7_c_RNI8D1A4_0_LC_9_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7498),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un61_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_RNILM0C_7_LC_9_9_6.C_ON=1'b0;
    defparam visibleX_RNILM0C_7_LC_9_9_6.SEQ_MODE=4'b0000;
    defparam visibleX_RNILM0C_7_LC_9_9_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 visibleX_RNILM0C_7_LC_9_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7489),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un54_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_9_LC_9_10_1.C_ON=1'b0;
    defparam visibleX_9_LC_9_10_1.SEQ_MODE=4'b1000;
    defparam visibleX_9_LC_9_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 visibleX_9_LC_9_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7468),
            .lcout(visibleXZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__7374),
            .ce(N__7298),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_9_11_0.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_9_11_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_9_11_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_LC_9_11_0 (
            .in0(_gnd_net_),
            .in1(N__7800),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8P8_LC_9_11_1.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8P8_LC_9_11_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8P8_LC_9_11_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8P8_LC_9_11_1 (
            .in0(_gnd_net_),
            .in1(N__7736),
            .in2(_gnd_net_),
            .in3(N__7243),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4_c_RNIV8PZ0Z8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_4),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQ8_LC_9_11_2.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQ8_LC_9_11_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQ8_LC_9_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQ8_LC_9_11_2 (
            .in0(_gnd_net_),
            .in1(N__7740),
            .in2(N__7769),
            .in3(N__7231),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5_c_RNI0BQZ0Z8),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_5),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_11_3.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_11_3.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_LUT4_0_LC_9_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7222),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6_THRU_CO),
            .ltout(),
            .carryin(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_6),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_11_4.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_11_4.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_LUT4_0_LC_9_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7219),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_cry_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam visibleX_RNINO0C_9_LC_9_11_7.C_ON=1'b0;
    defparam visibleX_RNINO0C_9_LC_9_11_7.SEQ_MODE=4'b0000;
    defparam visibleX_RNINO0C_9_LC_9_11_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 visibleX_RNINO0C_9_LC_9_11_7 (
            .in0(N__7801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_12_0.C_ON=1'b1;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_12_0.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_LC_9_12_0 (
            .in0(_gnd_net_),
            .in1(N__7770),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_LC_9_12_1.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_LC_9_12_1.LUT_INIT=16'b0000111111110000;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_LC_9_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7591),
            .in3(N__7582),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0),
            .ltout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGBZ0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_0_LC_9_12_2.C_ON=1'b0;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_0_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_0_LC_9_12_2.LUT_INIT=16'b0000111100001111;
    LogicCell40 chessboardpixel_un5_pixel_if_generate_plus_mult1_un33_sum_cry_6_c_RNI5JGB_0_LC_9_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7570),
            .in3(_gnd_net_),
            .lcout(chessboardpixel_un5_pixel_if_generate_plus_mult1_un40_sum_i_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam N_75_i_i_LC_12_16_1.C_ON=1'b0;
    defparam N_75_i_i_LC_12_16_1.SEQ_MODE=4'b0000;
    defparam N_75_i_i_LC_12_16_1.LUT_INIT=16'b1010101010011001;
    LogicCell40 N_75_i_i_LC_12_16_1 (
            .in0(N__7555),
            .in1(N__7509),
            .in2(_gnd_net_),
            .in3(N__7521),
            .lcout(G_256),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam N_555_i_LC_12_16_5.C_ON=1'b0;
    defparam N_555_i_LC_12_16_5.SEQ_MODE=4'b0000;
    defparam N_555_i_LC_12_16_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 N_555_i_LC_12_16_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7520),
            .lcout(G_255),
            .ltout(G_255_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CharacterDisplay.Z_decfrac15_0_a2_LC_12_16_6 .C_ON=1'b0;
    defparam \CharacterDisplay.Z_decfrac15_0_a2_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \CharacterDisplay.Z_decfrac15_0_a2_LC_12_16_6 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \CharacterDisplay.Z_decfrac15_0_a2_LC_12_16_6  (
            .in0(N__7508),
            .in1(_gnd_net_),
            .in2(N__7558),
            .in3(N__7554),
            .lcout(CharacterDisplay__decfrac8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SUM1_3_0_x2_LC_12_16_7.C_ON=1'b0;
    defparam SUM1_3_0_x2_LC_12_16_7.SEQ_MODE=4'b0000;
    defparam SUM1_3_0_x2_LC_12_16_7.LUT_INIT=16'b1100110000110011;
    LogicCell40 SUM1_3_0_x2_LC_12_16_7 (
            .in0(_gnd_net_),
            .in1(N__7510),
            .in2(_gnd_net_),
            .in3(N__7522),
            .lcout(G_254),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // SimpleVGA
